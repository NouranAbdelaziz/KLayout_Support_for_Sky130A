* Extracted by KLayout on : 15/07/2021 16:08

.SUBCKT mprj_logic_high
X$1 \$1 \$1 \$144 VNB sky130_fd_sc_hd__decap_6
X$2 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_3
X$3 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$4 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$5 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$6 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$7 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$8 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$9 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$10 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$11 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$12 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$13 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$14 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$15 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$16 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$17 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$18 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$20 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$21 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$22 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$23 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$24 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$25 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$26 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$27 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$28 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$29 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$30 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$31 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$32 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$33 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$34 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$35 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$36 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$37 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$40 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$41 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$42 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$43 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$44 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$45 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$46 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$47 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$48 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$49 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$50 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$51 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$52 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$53 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$54 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$55 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$56 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$57 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$60 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$61 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$62 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$63 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$64 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$65 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$66 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$67 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$68 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$69 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$70 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$71 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$72 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$73 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$74 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$75 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$76 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$77 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$80 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$81 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$82 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$83 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$84 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$85 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$86 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$87 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$88 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$89 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$90 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$91 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$92 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$93 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$94 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$95 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$96 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$97 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$100 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$101 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$102 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$103 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$104 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$105 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$106 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$107 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$108 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$109 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$110 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$111 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$112 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$113 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$114 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$115 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$116 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$117 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$120 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$121 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$122 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$123 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$124 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$125 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$126 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$127 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$128 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$131 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$132 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$133 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$134 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$135 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$136 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$137 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$138 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$139 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$140 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$141 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$142 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$143 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$144 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$145 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$146 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$147 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$148 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$151 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$152 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$153 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$154 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$155 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$156 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$157 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$158 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$159 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$160 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$161 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$162 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$163 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$164 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$165 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$166 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$167 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$168 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$171 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$172 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$173 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$174 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$175 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$176 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$177 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$178 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$179 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$180 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$181 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$182 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$183 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$184 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$185 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$186 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$187 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$188 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$191 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$192 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$193 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$194 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$195 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$196 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$197 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$198 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$199 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$200 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$201 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$202 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$203 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$204 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$205 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$206 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$207 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$208 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$211 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$212 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$213 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$214 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$215 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$216 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$217 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$218 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$219 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$220 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$221 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$222 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$223 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$224 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$225 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$226 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$227 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$228 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$231 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$232 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$233 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$234 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$235 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$236 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$237 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$238 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$239 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$240 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$241 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$242 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$243 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$244 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$245 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$246 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$247 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$248 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$251 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$252 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$253 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$254 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_8
X$255 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_3
X$256 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_3
X$257 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$258 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$259 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$260 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$261 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$264 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$265 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$266 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_4
X$268 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$269 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$270 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_4
X$272 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$273 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$274 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_4
X$276 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$277 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$278 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_4
X$280 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$281 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$282 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_4
X$284 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$285 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$286 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_4
X$288 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$289 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$290 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_4
X$292 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$293 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$294 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_4
X$296 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$297 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$298 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_4
X$300 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$301 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$302 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_4
X$304 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$305 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$306 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_4
X$308 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$309 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$310 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_4
X$312 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$313 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$314 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_4
X$316 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$317 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$318 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_4
X$320 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$321 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$322 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_4
X$324 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$325 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$326 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_4
X$328 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$329 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$330 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_4
X$332 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$333 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$334 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_4
X$336 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$337 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$338 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_4
X$340 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$341 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$342 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_4
X$344 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$345 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$346 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_4
X$348 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$349 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$350 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_4
X$352 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$353 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$354 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_4
X$356 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$357 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$358 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_4
X$360 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$361 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$362 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_4
X$364 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$365 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_8
X$367 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_3
X$368 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_3
X$369 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_3
X$370 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$371 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$372 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$373 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$374 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$375 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$376 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$379 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$380 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$381 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$383 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$384 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$385 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$386 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$387 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$388 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$390 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$391 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$392 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$393 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$394 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$395 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$396 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$397 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$398 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$401 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$402 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$403 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$405 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$406 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$407 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$409 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$410 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$413 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$414 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$415 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$416 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$417 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$419 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$421 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$422 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$425 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$427 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$428 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$429 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$430 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$431 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$432 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$433 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$434 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$437 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$438 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$440 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$441 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$442 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$443 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$444 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$445 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$448 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$449 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$451 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$452 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$453 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$454 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$455 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$456 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$459 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$460 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$461 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$462 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$464 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$465 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$466 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$467 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$468 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$470 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$471 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$472 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$473 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$474 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$475 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$477 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$479 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$482 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$483 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$484 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$485 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$486 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$487 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$488 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$489 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$490 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$493 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$494 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$495 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$496 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$497 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$498 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$499 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$500 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$502 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$504 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$505 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$506 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$507 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_8
X$510 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$511 \$1 \$1 \$144 VNB sky130_fd_sc_hd__decap_6
X$513 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$514 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$515 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$518 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$519 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$520 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$521 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$522 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$523 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$524 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$525 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$526 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$529 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$531 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$532 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$533 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$534 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$535 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$536 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$537 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$541 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$543 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$544 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$545 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$546 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$547 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$548 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$549 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$552 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$554 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$555 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$556 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$557 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$558 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$559 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$560 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$561 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_3
X$563 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$564 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$565 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$566 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$567 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$568 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$570 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$571 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$572 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$575 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$576 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$577 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$578 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$579 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$581 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$582 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$583 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$587 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$588 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$589 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$590 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$592 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$593 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$594 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$595 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$598 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$599 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$600 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$602 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$603 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$604 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$605 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$606 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$607 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$609 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$610 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$611 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$612 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$613 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$614 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$615 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$616 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$617 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$620 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$621 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$622 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$623 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$624 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$626 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$627 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$629 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$632 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$634 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$635 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$636 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$637 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$638 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$639 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$640 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$641 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$643 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$644 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$645 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$647 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$648 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$649 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$651 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$652 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$655 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$656 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$657 \$1 \$1 \$144 VNB sky130_fd_sc_hd__decap_6
X$659 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_3
X$660 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_3
X$661 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_3
X$662 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_8
X$663 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$665 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$666 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$667 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$668 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$670 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$671 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$672 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$673 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_4
X$674 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$676 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_4
X$678 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$679 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$680 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$681 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$682 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_8
X$683 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$686 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$687 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$688 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$689 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_8
X$690 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_8
X$692 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$693 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_3
X$694 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$695 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$696 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$697 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_3
X$698 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$699 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$701 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_8
X$702 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$703 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$704 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_4
X$706 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$707 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$708 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_8
X$710 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$711 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$712 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$713 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_4
X$714 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$715 \$1 \$1 \$144 VNB sky130_fd_sc_hd__decap_6
X$716 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$719 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$720 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$721 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$722 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$723 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_8
X$725 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_8
X$726 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$727 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$728 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$729 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$730 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_4
X$731 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$733 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$734 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$735 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$736 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_8
X$737 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$739 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$740 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$741 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$743 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$744 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_4
X$745 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$747 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$748 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$749 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$750 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_8
X$751 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$753 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$754 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_4
X$755 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$756 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$757 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$758 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$761 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$762 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$763 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$764 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_8
X$765 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$767 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$768 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$769 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$770 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_8
X$771 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$773 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_4
X$775 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$776 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$777 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$778 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$779 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_8
X$781 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$782 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$783 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$784 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$785 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_8
X$786 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$789 \$1 \$1 \$144 VNB sky130_fd_sc_hd__decap_6
X$790 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$791 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$792 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$793 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_8
X$794 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$796 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$797 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_4
X$799 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$800 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$801 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$802 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$803 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_3
X$805 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$806 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$807 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_8
X$809 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_8
X$810 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$811 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$813 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$814 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$815 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$816 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_4
X$818 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$819 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$821 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_8
X$822 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$823 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$824 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$825 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_8
X$826 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$828 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$829 \$1 \$1 \$144 VNB sky130_fd_sc_hd__decap_6
X$830 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$832 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$833 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_8
X$834 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_3
X$835 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$837 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$838 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$839 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$840 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_8
X$841 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$843 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$844 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$845 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$846 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_8
X$847 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$849 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$850 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$851 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$852 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$853 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_8
X$854 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$856 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$857 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_4
X$858 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$860 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$861 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_8
X$862 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$866 \$1 \$1 \$144 VNB sky130_fd_sc_hd__conb_1
X$867 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$868 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$869 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_12
X$870 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_8
X$872 \$1 \$1 \$144 VNB sky130_fd_sc_hd__decap_6
X$873 \$1 \$1 \$144 VNB sky130_fd_sc_hd__decap_6
X$874 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_3
X$875 \$1 \$144 \$1 VNB sky130_fd_sc_hd__decap_3
.ENDS mprj_logic_high

.SUBCKT sky130_fd_sc_hd__decap_8 VPB VGND VPWR VNB
M$1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=2890000U W=870000U
+ AS=226200000000P AD=226200000000P PS=2260000U PD=2260000U
M$2 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 L=2890000U W=550000U
+ AS=143000000000P AD=143000000000P PS=1620000U PD=1620000U
.ENDS sky130_fd_sc_hd__decap_8

.SUBCKT sky130_fd_sc_hd__decap_4 VPB VGND VPWR VNB
M$1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=1050000U W=870000U
+ AS=226200000000P AD=226200000000P PS=2260000U PD=2260000U
M$2 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 L=1050000U W=550000U
+ AS=143000000000P AD=143000000000P PS=1620000U PD=1620000U
.ENDS sky130_fd_sc_hd__decap_4

.SUBCKT sky130_fd_sc_hd__conb_1 VPB HI|VPWR LO|VGND VNB
R$1 LO|VGND LO|VGND 0
R$2 HI|VPWR HI|VPWR 0
.ENDS sky130_fd_sc_hd__conb_1

.SUBCKT sky130_fd_sc_hd__decap_3 VPB VGND VPWR VNB
M$1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=590000U W=870000U
+ AS=226200000000P AD=226200000000P PS=2260000U PD=2260000U
M$2 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 L=590000U W=550000U
+ AS=143000000000P AD=143000000000P PS=1620000U PD=1620000U
.ENDS sky130_fd_sc_hd__decap_3

.SUBCKT sky130_fd_sc_hd__decap_6 VPB VPWR VGND VNB
M$1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=1970000U W=870000U
+ AS=226200000000P AD=226200000000P PS=2260000U PD=2260000U
M$2 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 L=1970000U W=550000U
+ AS=143000000000P AD=143000000000P PS=1620000U PD=1620000U
.ENDS sky130_fd_sc_hd__decap_6

.SUBCKT sky130_fd_sc_hd__decap_12 VPB VGND VPWR VNB
M$1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=4730000U W=870000U
+ AS=226200000000P AD=226200000000P PS=2260000U PD=2260000U
M$2 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 L=4730000U W=550000U
+ AS=143000000000P AD=143000000000P PS=1620000U PD=1620000U
.ENDS sky130_fd_sc_hd__decap_12
