* Extracted by KLayout on : 15/07/2021 16:00

.SUBCKT digital_pll
X$1 \$3 \$114 \$1 \$252 \$249 \$3 \$18 VNB sky130_fd_sc_hd__mux2_1
X$2 \$18 \$54 \$70 \$2 \$61 \$76 \$77 \$3 \$3 VNB sky130_fd_sc_hd__o221ai_2
X$3 \$3 \$2 \$61 \$3 \$78 \$18 VNB sky130_fd_sc_hd__nand2_2
X$4 \$3 \$3 \$206 \$3 \$227 \$18 VNB sky130_fd_sc_hd__einvp_1
X$5 \$3 \$114 \$267 \$274 \$263 \$3 \$18 VNB sky130_fd_sc_hd__mux2_1
X$6 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$8 \$3 \$263 \$285 \$280 \$3 \$18 VNB sky130_fd_sc_hd__einvp_2
X$9 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$11 \$3 \$256 \$261 \$227 \$3 \$18 VNB sky130_fd_sc_hd__einvp_2
X$12 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$13 \$3 \$170 \$246 \$275 \$3 \$18 VNB sky130_fd_sc_hd__or2_2
X$15 \$3 \$114 \$83 \$275 \$282 \$3 \$18 VNB sky130_fd_sc_hd__mux2_1
X$16 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$19 \$3 \$114 \$233 \$270 \$272 \$3 \$18 VNB sky130_fd_sc_hd__mux2_1
X$21 \$3 \$242 \$18 \$3 \$200 VNB sky130_fd_sc_hd__inv_2
X$23 \$3 \$182 \$257 \$283 \$3 \$18 VNB sky130_fd_sc_hd__or2_2
X$25 \$3 \$114 \$277 \$246 \$151 \$3 \$18 VNB sky130_fd_sc_hd__mux2_1
X$27 \$3 \$114 \$278 \$230 \$284 \$3 \$18 VNB sky130_fd_sc_hd__mux2_1
X$29 \$3 \$276 \$279 \$273 \$3 \$18 VNB sky130_fd_sc_hd__einvp_2
X$32 \$18 \$271 \$276 \$273 \$3 \$3 VNB sky130_fd_sc_hd__einvn_8
X$33 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$34 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$35 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$37 \$3 \$291 \$3 \$18 \$285 VNB sky130_fd_sc_hd__clkinv_1
X$39 \$3 \$288 \$286 \$291 \$3 \$18 VNB sky130_fd_sc_hd__einvp_2
X$41 \$3 \$280 \$3 \$18 \$226 VNB sky130_fd_sc_hd__clkbuf_2
X$43 \$3 \$264 \$286 \$18 \$3 VNB sky130_fd_sc_hd__clkbuf_1
X$46 \$3 \$182 \$297 \$18 \$3 VNB sky130_fd_sc_hd__buf_1
X$48 \$3 \$227 \$3 \$18 \$292 VNB sky130_fd_sc_hd__clkbuf_2
X$49 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$50 \$3 \$219 \$246 \$274 \$3 \$18 VNB sky130_fd_sc_hd__or2_2
X$52 \$3 \$214 \$193 \$222 \$3 \$18 VNB sky130_fd_sc_hd__or2_2
X$53 \$3 \$3 \$18 VNB sky130_fd_sc_hd__decap_6
X$54 \$18 \$287 \$293 \$289 \$3 \$3 VNB sky130_fd_sc_hd__einvn_4
X$56 \$3 \$165 \$3 \$18 \$287 VNB sky130_fd_sc_hd__clkbuf_2
X$58 \$3 \$304 \$3 \$18 \$294 VNB sky130_fd_sc_hd__clkbuf_2
X$59 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$61 \$3 \$222 \$18 \$3 \$202 VNB sky130_fd_sc_hd__inv_2
X$63 \$18 \$296 \$295 \$284 \$3 \$3 VNB sky130_fd_sc_hd__einvn_4
X$64 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$66 \$18 \$271 \$266 \$272 \$3 \$3 VNB sky130_fd_sc_hd__einvn_4
X$67 \$3 \$3 \$18 VNB sky130_fd_sc_hd__decap_6
X$68 \$3 \$290 \$3 \$18 \$239 VNB sky130_fd_sc_hd__clkbuf_2
X$70 \$3 \$239 \$232 \$18 \$3 VNB sky130_fd_sc_hd__clkbuf_1
X$72 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$73 \$3 \$236 \$3 \$18 \$234 VNB sky130_fd_sc_hd__clkinv_1
X$74 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$76 \$3 \$220 \$234 \$229 \$3 \$18 VNB sky130_fd_sc_hd__einvp_2
X$78 \$3 \$226 \$240 \$18 \$3 VNB sky130_fd_sc_hd__clkbuf_1
X$80 \$18 \$229 \$237 \$227 \$3 \$3 VNB sky130_fd_sc_hd__einvn_8
X$81 \$3 \$3 \$18 VNB sky130_fd_sc_hd__decap_6
X$82 \$3 \$183 \$193 \$170 \$221 \$3 \$18 \$241 VNB sky130_fd_sc_hd__o31a_2
X$83 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$85 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$86 \$3 \$136 \$242 \$193 \$183 \$18 \$3 \$231 VNB sky130_fd_sc_hd__or4_2
X$88 \$3 \$225 \$134 \$218 \$3 \$18 VNB sky130_fd_sc_hd__or2_2
X$89 \$3 \$3 \$18 VNB sky130_fd_sc_hd__decap_6
X$90 \$3 \$213 \$183 \$218 \$3 \$18 \$164 VNB sky130_fd_sc_hd__or3_2
X$92 \$3 \$214 \$213 \$212 \$3 \$18 VNB sky130_fd_sc_hd__or2_2
X$94 \$3 \$182 \$214 \$193 \$242 \$235 \$3 \$18 VNB sky130_fd_sc_hd__a31o_2
X$96 \$3 \$243 \$238 \$3 \$190 \$18 VNB sky130_fd_sc_hd__and2_2
X$99 \$3 \$136 \$164 \$3 \$238 \$18 VNB sky130_fd_sc_hd__nand2_2
X$101 \$18 \$239 \$228 \$224 \$3 \$3 VNB sky130_fd_sc_hd__einvn_4
X$102 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$103 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$104 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$105 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$106 \$18 \$226 \$236 \$245 \$3 \$3 VNB sky130_fd_sc_hd__einvn_4
X$108 \$3 \$245 \$240 \$236 \$3 \$18 VNB sky130_fd_sc_hd__einvp_2
X$111 \$3 \$249 \$250 \$251 \$3 \$18 VNB sky130_fd_sc_hd__einvp_2
X$113 \$3 \$147 \$122 \$18 \$3 VNB sky130_fd_sc_hd__clkbuf_1
X$115 \$3 \$246 \$212 \$182 \$18 \$3 \$199 VNB sky130_fd_sc_hd__o21a_2
X$117 \$3 \$193 \$18 \$3 \$213 VNB sky130_fd_sc_hd__inv_2
X$119 \$18 \$116 \$136 \$222 \$225 \$247 \$270 \$3 \$3 VNB
+ sky130_fd_sc_hd__o311a_2
X$120 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$121 \$3 \$3 \$18 VNB sky130_fd_sc_hd__decap_6
X$123 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$124 \$18 \$253 \$199 \$242 \$182 \$193 \$183 \$3 \$3 VNB
+ sky130_fd_sc_hd__o41a_2
X$126 \$3 \$182 \$257 \$164 \$243 \$3 \$18 VNB sky130_fd_sc_hd__mux2_1
X$127 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$128 \$18 \$239 \$248 \$254 \$3 \$3 VNB sky130_fd_sc_hd__einvn_8
X$130 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$131 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$132 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$134 \$18 \$264 \$291 \$288 \$3 \$3 VNB sky130_fd_sc_hd__einvn_4
X$135 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$137 \$18 \$292 \$298 \$172 \$3 \$3 VNB sky130_fd_sc_hd__einvn_8
X$139 \$3 \$114 \$302 \$269 \$303 \$3 \$18 VNB sky130_fd_sc_hd__mux2_1
X$140 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$142 \$3 \$303 \$320 \$304 \$3 \$18 VNB sky130_fd_sc_hd__einvp_2
X$143 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$145 \$18 \$294 \$282 \$290 \$3 \$3 VNB sky130_fd_sc_hd__einvn_8
X$146 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$147 \$3 \$299 \$300 \$305 \$3 \$18 VNB sky130_fd_sc_hd__einvp_2
X$149 \$3 \$284 \$301 \$295 \$3 \$18 VNB sky130_fd_sc_hd__einvp_2
X$151 \$3 \$266 \$3 \$18 \$279 VNB sky130_fd_sc_hd__clkinv_1
X$154 \$3 \$273 \$3 \$18 \$296 VNB sky130_fd_sc_hd__clkbuf_2
X$156 \$3 \$271 \$268 \$18 \$3 VNB sky130_fd_sc_hd__clkbuf_1
X$157 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$159 \$3 \$228 \$3 \$18 \$259 VNB sky130_fd_sc_hd__clkinv_1
X$160 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$161 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$162 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$163 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$164 \$3 \$114 \$308 \$297 \$288 \$3 \$18 VNB sky130_fd_sc_hd__mux2_1
X$165 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$166 \$3 \$305 \$3 \$18 \$264 VNB sky130_fd_sc_hd__clkbuf_2
X$167 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$170 \$3 \$298 \$309 \$172 \$3 \$18 VNB sky130_fd_sc_hd__einvp_2
X$172 \$3 \$307 \$311 \$310 \$3 \$18 VNB sky130_fd_sc_hd__einvp_2
X$174 \$18 \$287 \$303 \$304 \$3 \$3 VNB sky130_fd_sc_hd__einvn_8
X$176 \$3 \$289 \$312 \$293 \$3 \$18 VNB sky130_fd_sc_hd__einvp_2
X$178 \$3 \$282 \$306 \$290 \$3 \$18 VNB sky130_fd_sc_hd__einvp_2
X$182 \$18 \$296 \$299 \$305 \$3 \$3 VNB sky130_fd_sc_hd__einvn_8
X$184 \$3 \$313 \$3 \$18 \$306 VNB sky130_fd_sc_hd__clkinv_1
X$186 \$3 \$296 \$301 \$18 \$3 VNB sky130_fd_sc_hd__clkbuf_1
X$187 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_12
X$188 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_8
X$189 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$190 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$191 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$192 \$3 \$114 \$258 \$221 \$245 \$3 \$18 VNB sky130_fd_sc_hd__mux2_1
X$194 \$3 \$206 \$256 \$237 \$3 \$18 VNB sky130_fd_sc_hd__or2_2
X$196 \$18 \$229 \$251 \$249 \$3 \$3 VNB sky130_fd_sc_hd__einvn_4
X$198 \$3 \$3 \$18 VNB sky130_fd_sc_hd__conb_1
X$200 \$3 \$182 \$214 \$193 \$170 \$260 \$3 \$18 VNB sky130_fd_sc_hd__a31o_2
X$202 \$3 \$251 \$3 \$18 \$261 VNB sky130_fd_sc_hd__clkinv_1
X$205 \$18 \$230 \$116 \$136 \$212 \$134 \$170 \$3 \$3 VNB
+ sky130_fd_sc_hd__o41a_2
X$206 \$3 \$3 \$18 VNB sky130_fd_sc_hd__decap_6
X$207 \$18 \$252 \$219 \$200 \$222 \$182 \$257 \$3 \$3 VNB
+ sky130_fd_sc_hd__o311a_2
X$208 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$210 \$3 \$242 \$212 \$182 \$246 \$3 \$18 \$255 VNB sky130_fd_sc_hd__o31a_2
X$212 \$3 \$242 \$222 \$257 \$3 \$18 VNB sky130_fd_sc_hd__or2_2
X$214 \$3 \$136 \$202 \$18 \$3 \$262 VNB sky130_fd_sc_hd__nor2_2
X$215 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$217 \$3 \$114 \$107 \$255 \$276 \$3 \$18 VNB sky130_fd_sc_hd__mux2_1
X$219 \$3 \$248 \$259 \$254 \$3 \$18 VNB sky130_fd_sc_hd__einvp_2
X$220 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$221 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$222 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$224 \$18 \$264 \$263 \$280 \$3 \$3 VNB sky130_fd_sc_hd__einvn_8
X$226 \$3 \$229 \$250 \$18 \$3 VNB sky130_fd_sc_hd__clkbuf_1
X$229 \$3 \$114 \$281 \$265 \$256 \$3 \$18 VNB sky130_fd_sc_hd__mux2_1
X$231 \$3 \$182 \$212 \$170 \$246 \$3 \$18 \$265 VNB sky130_fd_sc_hd__o31a_2
X$233 \$3 \$182 \$212 \$219 \$246 \$3 \$18 \$269 VNB sky130_fd_sc_hd__o31a_2
X$235 \$3 \$170 \$18 \$3 \$225 VNB sky130_fd_sc_hd__inv_2
X$237 \$18 \$270 \$170 \$134 \$222 \$182 \$257 \$3 \$3 VNB
+ sky130_fd_sc_hd__o311a_2
X$239 \$3 \$212 \$242 \$136 \$3 \$18 \$247 VNB sky130_fd_sc_hd__or3_2
X$240 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$243 \$3 \$114 \$15 \$262 \$289 \$3 \$18 VNB sky130_fd_sc_hd__mux2_1
X$245 \$3 \$182 \$222 \$246 \$3 \$18 VNB sky130_fd_sc_hd__or2_2
X$246 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$247 \$3 \$272 \$268 \$266 \$3 \$18 VNB sky130_fd_sc_hd__einvp_2
X$249 \$3 \$114 \$244 \$235 \$248 \$3 \$18 VNB sky130_fd_sc_hd__mux2_1
X$251 \$3 \$254 \$3 \$18 \$271 VNB sky130_fd_sc_hd__clkbuf_2
X$252 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$253 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$254 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$255 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$256 \$3 \$66 \$57 \$67 \$33 \$3 \$18 \$73 VNB sky130_fd_sc_hd__o211a_2
X$257 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$259 \$18 \$74 \$82 \$101 \$94 \$98 \$3 \$3 VNB sky130_fd_sc_hd__o2bb2a_2
X$260 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$261 \$18 \$46 \$82 \$5 \$84 \$3 \$3 VNB sky130_fd_sc_hd__dfrtp_2
X$262 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$264 \$3 \$77 \$76 \$25 \$87 \$18 \$51 \$3 VNB sky130_fd_sc_hd__a22o_2
X$265 \$3 \$3 \$18 VNB sky130_fd_sc_hd__decap_6
X$266 \$18 \$78 \$88 \$92 \$91 \$66 \$85 \$3 \$3 VNB sky130_fd_sc_hd__o221a_2
X$268 \$3 \$85 \$70 \$93 \$3 \$18 VNB sky130_fd_sc_hd__or2_2
X$269 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$270 \$18 \$86 \$55 \$5 \$95 \$3 \$3 VNB sky130_fd_sc_hd__dfrtp_2
X$273 \$3 \$32 \$55 \$52 \$24 \$18 \$95 \$3 VNB sky130_fd_sc_hd__a22o_2
X$275 \$3 \$60 \$18 \$3 \$72 VNB sky130_fd_sc_hd__inv_2
X$277 \$3 \$8 \$86 \$18 \$3 VNB sky130_fd_sc_hd__buf_1
X$278 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$279 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$280 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$281 \$3 \$57 \$18 \$3 \$91 VNB sky130_fd_sc_hd__inv_2
X$283 \$3 \$69 \$18 \$3 \$94 VNB sky130_fd_sc_hd__inv_2
X$285 \$3 \$82 \$101 \$18 \$3 \$98 VNB sky130_fd_sc_hd__nor2_2
X$287 \$3 \$82 \$98 \$101 \$3 \$75 \$18 VNB sky130_fd_sc_hd__a21oi_2
X$290 \$3 \$24 \$82 \$101 \$32 \$18 \$104 \$3 VNB sky130_fd_sc_hd__a22o_2
X$292 \$3 \$76 \$24 \$4 \$3 \$105 \$18 VNB sky130_fd_sc_hd__a21oi_2
X$293 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$295 \$3 \$24 \$25 \$87 \$32 \$18 \$99 \$3 VNB sky130_fd_sc_hd__a22o_2
X$297 \$3 \$25 \$18 \$3 \$76 VNB sky130_fd_sc_hd__inv_2
X$299 \$3 \$87 \$18 \$3 \$77 VNB sky130_fd_sc_hd__inv_2
X$300 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$301 \$3 \$73 \$18 \$3 \$88 VNB sky130_fd_sc_hd__inv_2
X$303 \$3 \$96 \$102 \$283 \$3 \$18 \$97 VNB sky130_fd_sc_hd__or3_2
X$306 \$18 \$62 \$93 \$97 \$71 \$70 \$106 \$3 \$3 VNB sky130_fd_sc_hd__o221a_2
X$308 \$3 \$44 \$79 \$43 \$3 \$92 \$18 VNB sky130_fd_sc_hd__a21oi_2
X$310 \$3 \$81 \$18 \$3 \$80 VNB sky130_fd_sc_hd__inv_2
X$311 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$312 \$18 \$130 \$108 \$5 \$100 \$3 \$3 VNB sky130_fd_sc_hd__dfrtp_2
X$314 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$316 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$317 \$3 \$8 \$103 \$18 \$3 VNB sky130_fd_sc_hd__buf_1
X$319 \$18 \$103 \$101 \$5 \$104 \$3 \$3 VNB sky130_fd_sc_hd__dfrtp_2
X$321 \$18 \$156 \$25 \$5 \$105 \$3 \$3 VNB sky130_fd_sc_hd__dfrtp_2
X$322 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$324 \$3 \$82 \$18 \$3 \$53 VNB sky130_fd_sc_hd__inv_2
X$325 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$326 \$18 \$140 \$96 \$5 \$110 \$3 \$3 VNB sky130_fd_sc_hd__dfrtp_2
X$327 \$3 \$3 \$18 VNB sky130_fd_sc_hd__decap_6
X$328 \$18 \$109 \$102 \$5 \$111 \$3 \$3 VNB sky130_fd_sc_hd__dfrtp_2
X$331 \$3 \$32 \$18 \$3 \$24 VNB sky130_fd_sc_hd__inv_2
X$332 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$334 \$18 \$32 \$100 \$100 \$108 \$108 \$3 \$3 VNB sky130_fd_sc_hd__a2bb2o_2
X$335 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$336 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$337 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$338 \$3 \$114 \$129 \$116 \$128 \$3 \$18 VNB sky130_fd_sc_hd__mux2_1
X$339 \$3 \$3 \$18 VNB sky130_fd_sc_hd__decap_6
X$340 \$3 \$117 \$205 \$115 \$3 \$18 VNB sky130_fd_sc_hd__einvp_2
X$341 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$344 \$3 \$118 \$122 \$119 \$3 \$18 VNB sky130_fd_sc_hd__einvp_2
X$345 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$347 \$3 \$112 \$18 \$3 \$113 VNB sky130_fd_sc_hd__inv_2
X$349 \$18 \$168 \$87 \$5 \$99 \$3 \$3 VNB sky130_fd_sc_hd__dfrtp_2
X$350 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$351 \$3 \$120 \$113 \$112 \$96 \$3 \$110 \$18 VNB sky130_fd_sc_hd__o22a_2
X$352 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$354 \$3 \$102 \$18 \$3 \$124 VNB sky130_fd_sc_hd__inv_2
X$356 \$18 \$113 \$111 \$121 \$112 \$124 \$3 \$3 VNB sky130_fd_sc_hd__o22ai_2
X$357 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$358 \$3 \$125 \$3 \$18 \$147 VNB sky130_fd_sc_hd__clkbuf_2
X$360 \$18 \$127 \$100 \$5 \$126 \$3 \$3 VNB sky130_fd_sc_hd__dfrtp_2
X$361 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$362 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$363 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$364 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$366 \$18 \$67 \$33 \$66 \$56 \$50 \$3 \$3 VNB sky130_fd_sc_hd__a22oi_2
X$367 \$3 \$56 \$50 \$57 \$3 \$18 VNB sky130_fd_sc_hd__or2_2
X$369 \$18 \$8 \$40 \$5 \$39 \$3 \$3 VNB sky130_fd_sc_hd__dfrtp_2
X$371 \$18 \$50 \$68 \$68 \$74 \$74 \$3 \$3 VNB sky130_fd_sc_hd__a2bb2o_2
X$372 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$375 \$18 \$67 \$69 \$69 \$75 \$75 \$3 \$3 VNB sky130_fd_sc_hd__a2bb2o_2
X$377 \$18 \$58 \$30 \$40 \$74 \$38 \$3 \$3 VNB sky130_fd_sc_hd__o2bb2a_2
X$378 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$380 \$3 \$47 \$32 \$10 \$59 \$84 \$3 \$18 VNB sky130_fd_sc_hd__a31o_2
X$382 \$3 \$34 \$28 \$53 \$18 \$59 \$3 VNB sky130_fd_sc_hd__o21ai_2
X$384 \$3 \$28 \$34 \$53 \$3 \$18 \$10 VNB sky130_fd_sc_hd__or3_2
X$385 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$388 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$389 \$3 \$54 \$51 \$58 \$3 \$18 \$61 VNB sky130_fd_sc_hd__a21bo_2
X$391 \$3 \$51 \$58 \$54 \$3 \$18 VNB sky130_fd_sc_hd__or2_2
X$394 \$3 \$47 \$48 \$29 \$3 \$18 VNB sky130_fd_sc_hd__or2_2
X$396 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$397 \$3 \$28 \$37 \$41 \$3 \$60 \$18 VNB sky130_fd_sc_hd__a21oi_2
X$399 \$18 \$78 \$71 \$73 \$79 \$60 \$80 \$3 \$3 VNB sky130_fd_sc_hd__o2111ai_2
X$401 \$3 \$42 \$37 \$26 \$20 \$18 \$69 \$3 VNB sky130_fd_sc_hd__a22o_2
X$403 \$18 \$45 \$81 \$72 \$43 \$44 \$79 \$3 \$3 VNB sky130_fd_sc_hd__o221a_2
X$404 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$405 \$3 \$49 \$55 \$24 \$52 \$3 \$18 \$62 VNB sky130_fd_sc_hd__and4_2
X$406 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$408 \$18 \$64 \$52 \$5 \$63 \$3 \$3 VNB sky130_fd_sc_hd__dfrtp_2
X$410 \$3 \$24 \$49 \$52 \$32 \$18 \$63 \$3 VNB sky130_fd_sc_hd__a22o_2
X$412 \$3 \$8 \$64 \$18 \$3 VNB sky130_fd_sc_hd__buf_1
X$414 \$3 \$143 \$65 \$18 \$3 VNB sky130_fd_sc_hd__clkbuf_1
X$415 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$417 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$418 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$419 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$420 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$421 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$422 \$3 \$3 \$18 VNB sky130_fd_sc_hd__decap_6
X$424 \$3 \$8 \$46 \$18 \$3 VNB sky130_fd_sc_hd__buf_1
X$426 \$18 \$17 \$30 \$5 \$23 \$3 \$3 VNB sky130_fd_sc_hd__dfrtp_2
X$428 \$3 \$30 \$40 \$18 \$3 \$38 VNB sky130_fd_sc_hd__nor2_2
X$430 \$3 \$38 \$30 \$40 \$3 \$18 \$68 VNB sky130_fd_sc_hd__a21o_2
X$433 \$3 \$24 \$30 \$40 \$32 \$18 \$39 \$3 VNB sky130_fd_sc_hd__a22o_2
X$434 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$435 \$18 \$32 \$25 \$4 \$9 \$30 \$23 \$3 \$3 VNB sky130_fd_sc_hd__o221a_2
X$436 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$437 \$3 \$32 \$25 \$9 \$30 \$3 \$18 \$47 VNB sky130_fd_sc_hd__and4_2
X$439 \$18 \$6 \$25 \$9 \$30 \$28 \$24 \$3 \$3 VNB sky130_fd_sc_hd__a311o_2
X$441 \$3 \$5 \$18 \$36 \$3 VNB sky130_fd_sc_hd__buf_2
X$445 \$18 \$32 \$26 \$12 \$28 \$34 \$48 \$3 \$3 VNB sky130_fd_sc_hd__o221a_2
X$447 \$3 \$26 \$18 \$3 \$34 VNB sky130_fd_sc_hd__inv_2
X$449 \$18 \$22 \$26 \$5 \$29 \$3 \$3 VNB sky130_fd_sc_hd__dfrtp_2
X$451 \$3 \$24 \$12 \$19 \$32 \$18 \$13 \$3 VNB sky130_fd_sc_hd__a22o_2
X$453 \$3 \$28 \$41 \$18 \$3 \$37 VNB sky130_fd_sc_hd__nor2_2
X$458 \$3 \$19 \$18 \$3 \$41 VNB sky130_fd_sc_hd__inv_2
X$459 \$18 \$37 \$42 \$43 \$37 \$42 \$3 \$3 VNB sky130_fd_sc_hd__o2bb2ai_2
X$460 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$461 \$18 \$42 \$26 \$20 \$20 \$26 \$3 \$3 VNB sky130_fd_sc_hd__o2bb2a_2
X$463 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$464 \$3 \$44 \$43 \$3 \$45 \$18 VNB sky130_fd_sc_hd__nand2_2
X$465 \$3 \$49 \$24 \$31 \$3 \$18 VNB sky130_fd_sc_hd__or2_2
X$466 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$467 \$18 \$21 \$49 \$5 \$31 \$3 \$3 VNB sky130_fd_sc_hd__dfrtp_2
X$470 \$3 \$24 \$26 \$20 \$32 \$18 \$7 \$3 VNB sky130_fd_sc_hd__a22o_2
X$472 \$3 \$8 \$22 \$18 \$3 VNB sky130_fd_sc_hd__buf_1
X$474 \$3 \$27 \$3 \$18 \$35 VNB sky130_fd_sc_hd__clkinv_1
X$475 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$476 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$477 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$478 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$479 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_8
X$480 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$482 \$3 \$8 \$11 \$18 \$3 VNB sky130_fd_sc_hd__buf_1
X$484 \$3 \$8 \$17 \$18 \$3 VNB sky130_fd_sc_hd__buf_1
X$486 \$3 \$30 \$9 \$3 \$4 \$18 VNB sky130_fd_sc_hd__nand2_2
X$489 \$3 \$10 \$18 \$3 \$9 VNB sky130_fd_sc_hd__inv_2
X$491 \$18 \$11 \$12 \$5 \$6 \$3 \$3 VNB sky130_fd_sc_hd__dfrtp_2
X$494 \$3 \$12 \$18 \$3 \$28 VNB sky130_fd_sc_hd__inv_2
X$496 \$18 \$14 \$19 \$5 \$13 \$3 \$3 VNB sky130_fd_sc_hd__dfrtp_2
X$499 \$3 \$8 \$14 \$18 \$3 VNB sky130_fd_sc_hd__buf_1
X$501 \$18 \$16 \$20 \$5 \$7 \$3 \$3 VNB sky130_fd_sc_hd__dfrtp_2
X$504 \$3 \$8 \$16 \$18 \$3 VNB sky130_fd_sc_hd__buf_1
X$506 \$3 \$8 \$21 \$18 \$3 VNB sky130_fd_sc_hd__buf_1
X$507 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_8
X$508 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$509 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$510 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$511 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$514 \$3 \$132 \$138 \$18 \$3 VNB sky130_fd_sc_hd__clkbuf_1
X$515 \$18 \$167 \$162 \$159 \$3 \$3 VNB sky130_fd_sc_hd__einvn_8
X$517 \$3 \$162 \$163 \$159 \$3 \$18 VNB sky130_fd_sc_hd__einvp_2
X$519 \$3 \$159 \$3 \$18 \$132 VNB sky130_fd_sc_hd__clkbuf_2
X$521 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$522 \$3 \$8 \$168 \$18 \$3 VNB sky130_fd_sc_hd__buf_1
X$523 \$3 \$8 \$156 \$18 \$3 VNB sky130_fd_sc_hd__buf_1
X$527 \$3 \$172 \$3 \$18 \$167 VNB sky130_fd_sc_hd__clkbuf_2
X$528 \$18 \$147 \$119 \$118 \$3 \$3 VNB sky130_fd_sc_hd__einvn_4
X$529 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$530 \$18 \$178 \$170 \$169 \$169 \$170 \$3 \$3 VNB sky130_fd_sc_hd__o2bb2a_2
X$531 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$532 \$3 \$150 \$195 \$165 \$3 \$18 VNB sky130_fd_sc_hd__einvp_2
X$534 \$3 \$8 \$179 \$18 \$3 VNB sky130_fd_sc_hd__buf_1
X$535 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$536 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$537 \$3 \$114 \$171 \$180 \$187 \$3 \$18 VNB sky130_fd_sc_hd__mux2_1
X$540 \$3 \$114 \$157 \$160 \$150 \$3 \$18 VNB sky130_fd_sc_hd__mux2_1
X$542 \$3 \$144 \$18 \$3 \$134 VNB sky130_fd_sc_hd__inv_2
X$543 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$545 \$18 \$148 \$113 \$149 \$144 \$112 \$145 \$3 \$3 VNB
+ sky130_fd_sc_hd__a32o_2
X$546 \$3 \$133 \$131 \$144 \$135 \$3 \$18 VNB sky130_fd_sc_hd__mux2_1
X$547 \$3 \$3 \$18 VNB sky130_fd_sc_hd__decap_6
X$548 \$3 \$3 \$18 VNB sky130_fd_sc_hd__decap_6
X$549 \$3 \$120 \$137 \$93 \$124 \$3 \$133 \$18 VNB sky130_fd_sc_hd__o22a_2
X$551 \$18 \$113 \$166 \$173 \$174 \$158 \$181 \$3 \$3 VNB
+ sky130_fd_sc_hd__a221o_2
X$553 \$3 \$120 \$124 \$164 \$3 \$18 \$142 VNB sky130_fd_sc_hd__or3_2
X$554 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$555 \$18 \$176 \$182 \$5 \$175 \$3 \$3 VNB sky130_fd_sc_hd__dfrtp_2
X$556 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$557 \$3 \$151 \$35 \$125 \$3 \$18 VNB sky130_fd_sc_hd__einvp_2
X$560 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$561 \$3 \$161 \$65 \$27 \$3 \$18 VNB sky130_fd_sc_hd__einvp_2
X$563 \$18 \$143 \$27 \$161 \$3 \$3 VNB sky130_fd_sc_hd__einvn_4
X$565 \$3 \$158 \$18 \$3 \$166 VNB sky130_fd_sc_hd__inv_2
X$566 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$567 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$569 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$570 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$571 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$572 \$3 \$128 \$138 \$139 \$3 \$18 VNB sky130_fd_sc_hd__einvp_2
X$574 \$18 \$132 \$117 \$115 \$3 \$3 VNB sky130_fd_sc_hd__einvn_8
X$575 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$577 \$3 \$8 \$140 \$18 \$3 VNB sky130_fd_sc_hd__buf_1
X$579 \$3 \$114 \$141 \$199 \$117 \$3 \$18 VNB sky130_fd_sc_hd__mux2_1
X$580 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$581 \$3 \$93 \$18 \$3 \$131 VNB sky130_fd_sc_hd__inv_2
X$584 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$585 \$3 \$133 \$123 \$3 \$145 \$18 VNB sky130_fd_sc_hd__nand2_2
X$587 \$3 \$135 \$112 \$93 \$134 \$3 \$18 \$169 VNB sky130_fd_sc_hd__o211a_2
X$588 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$590 \$3 \$136 \$131 \$142 \$106 \$3 \$18 \$112 VNB sky130_fd_sc_hd__o31a_2
X$592 \$18 \$121 \$120 \$120 \$137 \$137 \$3 \$3 VNB sky130_fd_sc_hd__a2bb2o_2
X$594 \$3 \$93 \$124 \$102 \$131 \$18 \$137 \$3 VNB sky130_fd_sc_hd__a22o_2
X$595 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$597 \$3 \$115 \$3 \$18 \$143 VNB sky130_fd_sc_hd__clkbuf_2
X$599 \$3 \$8 \$109 \$18 \$3 VNB sky130_fd_sc_hd__buf_1
X$601 \$3 \$8 \$130 \$18 \$3 VNB sky130_fd_sc_hd__buf_1
X$603 \$3 \$8 \$127 \$18 \$3 VNB sky130_fd_sc_hd__buf_1
X$605 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$606 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$608 \$18 \$132 \$139 \$128 \$3 \$3 VNB sky130_fd_sc_hd__einvn_4
X$610 \$3 \$114 \$153 \$154 \$118 \$3 \$18 VNB sky130_fd_sc_hd__mux2_1
X$613 \$3 \$8 \$146 \$18 \$3 VNB sky130_fd_sc_hd__buf_1
X$615 \$18 \$147 \$150 \$165 \$3 \$3 VNB sky130_fd_sc_hd__einvn_8
X$617 \$18 \$146 \$144 \$5 \$148 \$3 \$3 VNB sky130_fd_sc_hd__dfrtp_2
X$619 \$3 \$133 \$123 \$149 \$3 \$18 VNB sky130_fd_sc_hd__or2_2
X$620 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$622 \$3 \$96 \$18 \$3 \$120 VNB sky130_fd_sc_hd__inv_2
X$623 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$624 \$18 \$143 \$151 \$125 \$3 \$3 VNB sky130_fd_sc_hd__einvn_8
X$626 \$18 \$155 \$126 \$5 \$152 \$3 \$3 VNB sky130_fd_sc_hd__dfrtp_2
X$628 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$629 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$630 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$631 \$18 \$226 \$220 \$229 \$3 \$3 VNB sky130_fd_sc_hd__einvn_8
X$632 \$3 \$114 \$90 \$215 \$220 \$3 \$18 VNB sky130_fd_sc_hd__mux2_1
X$633 \$3 \$3 \$18 VNB sky130_fd_sc_hd__decap_6
X$634 \$3 \$186 \$3 \$18 \$163 VNB sky130_fd_sc_hd__clkinv_1
X$637 \$3 \$227 \$217 \$3 \$18 VNB sky130_fd_sc_hd__clkinv_2
X$638 \$3 \$216 \$89 \$3 \$206 \$18 VNB sky130_fd_sc_hd__nand2_2
X$640 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$642 \$3 \$114 \$206 \$18 \$3 \$8 VNB sky130_fd_sc_hd__nor2_2
X$643 \$18 \$5 \$217 \$3 \$3 VNB sky130_fd_sc_hd__clkinv_8
X$644 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$646 \$18 \$215 \$199 \$219 \$182 \$193 \$183 \$3 \$3 VNB
+ sky130_fd_sc_hd__o41a_2
X$647 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$648 \$3 \$182 \$222 \$212 \$18 \$3 \$221 VNB sky130_fd_sc_hd__and3_2
X$649 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$650 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$652 \$18 \$154 \$230 \$212 \$136 \$144 \$225 \$3 \$3 VNB
+ sky130_fd_sc_hd__o41a_2
X$655 \$3 \$218 \$18 \$3 \$219 VNB sky130_fd_sc_hd__inv_2
X$657 \$3 \$170 \$144 \$242 \$3 \$18 VNB sky130_fd_sc_hd__or2_2
X$659 \$18 \$180 \$136 \$212 \$225 \$231 \$230 \$3 \$3 VNB
+ sky130_fd_sc_hd__o311a_2
X$660 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$661 \$18 \$207 \$113 \$192 \$193 \$112 \$194 \$3 \$3 VNB
+ sky130_fd_sc_hd__a32o_2
X$663 \$3 \$219 \$200 \$18 \$3 \$201 VNB sky130_fd_sc_hd__nor2_2
X$665 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$666 \$3 \$93 \$213 \$193 \$131 \$18 \$189 \$3 VNB sky130_fd_sc_hd__a22o_2
X$668 \$3 \$213 \$93 \$192 \$18 \$204 \$3 VNB sky130_fd_sc_hd__o21ai_2
X$670 \$3 \$214 \$93 \$131 \$183 \$3 \$203 \$18 VNB sky130_fd_sc_hd__o22a_2
X$672 \$3 \$182 \$18 \$3 \$136 VNB sky130_fd_sc_hd__inv_2
X$674 \$18 \$210 \$214 \$5 \$223 \$3 \$3 VNB sky130_fd_sc_hd__dfrtp_2
X$676 \$3 \$183 \$112 \$209 \$18 \$223 \$3 VNB sky130_fd_sc_hd__o21ai_2
X$677 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$679 \$3 \$214 \$18 \$3 \$183 VNB sky130_fd_sc_hd__inv_2
X$680 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$681 \$3 \$114 \$211 \$241 \$224 \$3 \$18 VNB sky130_fd_sc_hd__mux2_1
X$683 \$3 \$224 \$232 \$228 \$3 \$18 VNB sky130_fd_sc_hd__einvp_2
X$684 \$3 \$3 \$18 VNB sky130_fd_sc_hd__decap_6
X$685 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$687 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$688 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$689 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$690 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$691 \$3 \$114 \$177 \$185 \$162 \$3 \$18 VNB sky130_fd_sc_hd__mux2_1
X$692 \$3 \$119 \$3 \$18 \$195 VNB sky130_fd_sc_hd__clkinv_1
X$694 \$3 \$139 \$3 \$18 \$205 VNB sky130_fd_sc_hd__clkinv_1
X$697 \$3 \$167 \$196 \$18 \$3 VNB sky130_fd_sc_hd__clkbuf_1
X$698 \$18 \$167 \$186 \$187 \$3 \$3 VNB sky130_fd_sc_hd__einvn_4
X$700 \$3 \$187 \$196 \$186 \$3 \$18 VNB sky130_fd_sc_hd__einvp_2
X$702 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$703 \$18 \$179 \$170 \$5 \$178 \$3 \$3 VNB sky130_fd_sc_hd__dfrtp_2
X$705 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$706 \$3 \$183 \$193 \$182 \$199 \$3 \$18 \$185 VNB sky130_fd_sc_hd__o31a_2
X$708 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$709 \$18 \$191 \$193 \$5 \$207 \$3 \$3 VNB sky130_fd_sc_hd__dfrtp_2
X$710 \$3 \$8 \$191 \$18 \$3 VNB sky130_fd_sc_hd__buf_1
X$713 \$18 \$160 \$199 \$170 \$182 \$193 \$183 \$3 \$3 VNB
+ sky130_fd_sc_hd__o41a_2
X$714 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$715 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$716 \$3 \$93 \$134 \$144 \$131 \$18 \$123 \$3 VNB sky130_fd_sc_hd__a22o_2
X$717 \$18 \$188 \$201 \$123 \$133 \$200 \$93 \$3 \$3 VNB
+ sky130_fd_sc_hd__o32a_2
X$719 \$3 \$188 \$189 \$192 \$3 \$18 VNB sky130_fd_sc_hd__or2_2
X$720 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$723 \$18 \$173 \$189 \$203 \$188 \$202 \$93 \$3 \$3 VNB
+ sky130_fd_sc_hd__o32a_2
X$724 \$3 \$136 \$93 \$131 \$182 \$3 \$158 \$18 VNB sky130_fd_sc_hd__o22a_2
X$727 \$3 \$136 \$112 \$181 \$18 \$175 \$3 VNB sky130_fd_sc_hd__o21ai_2
X$728 \$18 \$113 \$197 \$203 \$208 \$204 \$209 \$3 \$3 VNB
+ sky130_fd_sc_hd__a221o_2
X$731 \$3 \$173 \$18 \$3 \$174 VNB sky130_fd_sc_hd__inv_2
X$732 \$3 \$188 \$189 \$3 \$194 \$18 VNB sky130_fd_sc_hd__nand2_2
X$733 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$736 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$737 \$3 \$203 \$18 \$3 \$208 VNB sky130_fd_sc_hd__inv_2
X$739 \$3 \$114 \$184 \$190 \$161 \$3 \$18 VNB sky130_fd_sc_hd__mux2_1
X$740 \$3 \$204 \$18 \$3 \$197 VNB sky130_fd_sc_hd__inv_2
X$742 \$3 \$8 \$210 \$18 \$3 VNB sky130_fd_sc_hd__buf_1
X$745 \$3 \$8 \$176 \$18 \$3 VNB sky130_fd_sc_hd__buf_1
X$746 \$3 \$8 \$155 \$18 \$3 VNB sky130_fd_sc_hd__buf_1
X$747 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$749 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$750 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$751 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$752 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$753 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_12
X$754 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_12
X$755 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_12
X$756 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_12
X$759 \$18 \$292 \$310 \$307 \$3 \$3 VNB sky130_fd_sc_hd__einvn_4
X$762 \$3 \$310 \$3 \$18 \$309 VNB sky130_fd_sc_hd__clkinv_1
X$764 \$3 \$114 \$322 \$260 \$307 \$3 \$18 VNB sky130_fd_sc_hd__mux2_1
X$766 \$18 \$319 \$314 \$3 \$3 VNB sky130_fd_sc_hd__clkinv_8
X$768 \$3 \$292 \$311 \$18 \$3 VNB sky130_fd_sc_hd__clkbuf_1
X$769 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$770 \$3 \$293 \$3 \$18 \$320 VNB sky130_fd_sc_hd__clkinv_1
X$774 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$776 \$3 \$304 \$314 \$3 \$18 VNB sky130_fd_sc_hd__clkinv_2
X$777 \$3 \$114 \$317 \$283 \$298 \$3 \$18 VNB sky130_fd_sc_hd__mux2_1
X$778 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$779 \$3 \$287 \$312 \$18 \$3 VNB sky130_fd_sc_hd__clkbuf_1
X$780 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$781 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$782 \$18 \$294 \$313 \$315 \$3 \$3 VNB sky130_fd_sc_hd__einvn_4
X$784 \$3 \$315 \$321 \$313 \$3 \$18 VNB sky130_fd_sc_hd__einvp_2
X$785 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$786 \$3 \$3 \$18 VNB sky130_fd_sc_hd__decap_6
X$789 \$3 \$294 \$321 \$18 \$3 VNB sky130_fd_sc_hd__clkbuf_1
X$790 \$3 \$114 \$318 \$253 \$299 \$3 \$18 VNB sky130_fd_sc_hd__mux2_1
X$791 \$3 \$3 \$18 VNB sky130_fd_sc_hd__decap_6
X$792 \$3 \$295 \$3 \$18 \$300 VNB sky130_fd_sc_hd__clkinv_1
X$793 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$794 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_12
X$795 \$3 \$114 \$316 \$238 \$315 \$3 \$18 VNB sky130_fd_sc_hd__mux2_1
X$797 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_4
X$799 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_12
X$801 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_12
X$802 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_8
X$803 \$3 \$3 \$18 VNB sky130_fd_sc_hd__decap_6
X$806 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
X$807 \$3 \$18 \$3 VNB sky130_fd_sc_hd__decap_3
.ENDS digital_pll

.SUBCKT sky130_fd_sc_hd__o2bb2ai_2 VGND A1_N A2_N Y B1 B2 VPWR VPB VNB
M$1 VPWR A1_N \$6 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=280000000000P AD=135000000000P PS=2560000U PD=1270000U
M$2 \$6 A2_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$3 VPWR A2_N \$6 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$4 \$6 A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=400000000000P PS=1270000U PD=1800000U
M$5 VPWR \$6 Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=400000000000P AD=135000000000P PS=1800000U PD=1270000U
M$6 Y \$6 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=152500000000P PS=1270000U PD=1305000U
M$7 VPWR B1 \$12 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=152500000000P AD=135000000000P PS=1305000U PD=1270000U
M$8 \$12 B2 Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$9 Y B2 \$12 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$10 \$12 B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=285000000000P PS=1270000U PD=2570000U
M$11 \$7 \$6 Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=175500000000P
+ AD=87750000000P PS=1840000U PD=920000U
M$12 Y \$6 \$7 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=99125000000P PS=920000U PD=955000U
M$13 \$7 B1 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=99125000000P AD=87750000000P PS=955000U PD=920000U
M$14 VGND B2 \$7 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=87750000000P PS=920000U PD=920000U
M$15 \$7 B2 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=87750000000P PS=920000U PD=920000U
M$16 VGND B1 \$7 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=169000000000P PS=920000U PD=1820000U
M$17 VGND A1_N \$4 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=182000000000P AD=87750000000P PS=1860000U PD=920000U
M$18 \$4 A2_N \$6 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=87750000000P PS=920000U PD=920000U
M$19 \$6 A2_N \$4 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=87750000000P PS=920000U PD=920000U
M$20 \$4 A1_N VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=169000000000P PS=920000U PD=1820000U
.ENDS sky130_fd_sc_hd__o2bb2ai_2

.SUBCKT sky130_fd_sc_hd__o2111ai_2 VGND D1 Y C1 B1 A2 A1 VPWR VPB VNB
M$1 \$13 A2 Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=295000000000P AD=140000000000P PS=2590000U PD=1280000U
M$2 Y A2 \$13 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$3 \$13 A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$4 VPWR A1 \$13 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=330000000000P PS=1280000U PD=2660000U
M$5 VPWR D1 Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=265000000000P AD=140000000000P PS=2530000U PD=1280000U
M$6 Y D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$7 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$8 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$9 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$10 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=265000000000P PS=1280000U PD=2530000U
M$11 \$9 B1 \$7 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=175500000000P AD=91000000000P PS=1840000U PD=930000U
M$12 \$7 B1 \$9 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=91000000000P
+ AD=91000000000P PS=930000U PD=930000U
M$13 \$9 A2 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=91000000000P AD=91000000000P PS=930000U PD=930000U
M$14 VGND A2 \$9 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=91000000000P AD=91000000000P PS=930000U PD=930000U
M$15 \$9 A1 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=91000000000P AD=91000000000P PS=930000U PD=930000U
M$16 VGND A1 \$9 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=91000000000P AD=214500000000P PS=930000U PD=1960000U
M$17 \$4 D1 Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=224250000000P
+ AD=91000000000P PS=1990000U PD=930000U
M$18 Y D1 \$4 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=91000000000P
+ AD=91000000000P PS=930000U PD=930000U
M$19 \$4 C1 \$7 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=91000000000P
+ AD=91000000000P PS=930000U PD=930000U
M$20 \$7 C1 \$4 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=91000000000P
+ AD=191750000000P PS=930000U PD=1890000U
.ENDS sky130_fd_sc_hd__o2111ai_2

.SUBCKT sky130_fd_sc_hd__o22ai_2 VGND B1 Y B2 A2 A1 VPWR VPB VNB
M$1 \$11 A2 Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=280000000000P AD=135000000000P PS=2560000U PD=1270000U
M$2 Y A2 \$11 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$3 \$11 A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$4 VPWR A1 \$11 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=280000000000P PS=1270000U PD=2560000U
M$5 \$9 B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=280000000000P AD=135000000000P PS=2560000U PD=1270000U
M$6 VPWR B1 \$9 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$7 \$9 B2 Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$8 Y B2 \$9 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=280000000000P PS=1270000U PD=2560000U
M$9 \$3 B1 Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=182000000000P
+ AD=87750000000P PS=1860000U PD=920000U
M$10 Y B1 \$3 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$11 \$3 B2 Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$12 Y B2 \$3 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=269750000000P PS=920000U PD=1480000U
M$13 \$3 A2 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=269750000000P AD=87750000000P PS=1480000U PD=920000U
M$14 VGND A2 \$3 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=87750000000P PS=920000U PD=920000U
M$15 \$3 A1 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=87750000000P PS=920000U PD=920000U
M$16 VGND A1 \$3 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=169000000000P PS=920000U PD=1820000U
.ENDS sky130_fd_sc_hd__o22ai_2

.SUBCKT sky130_fd_sc_hd__a21bo_2 VPB B1_N A1 A2 VPWR VGND X VNB
M$1 \$11 \$10 \$6 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=135000000000P PS=2520000U PD=1270000U
M$2 \$6 A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$3 VPWR A2 \$6 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$4 \$10 B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=109200000000P AD=181500000000P PS=1360000U PD=1510000U
M$5 VPWR \$11 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=140000000000P PS=2520000U PD=1280000U
M$6 X \$11 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=181500000000P PS=1280000U PD=1510000U
M$7 VGND \$10 \$11 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=169000000000P AD=107250000000P PS=1820000U PD=980000U
M$8 \$11 A1 \$12 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=107250000000P AD=68250000000P PS=980000U PD=860000U
M$9 \$12 A2 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=68250000000P AD=169000000000P PS=860000U PD=1820000U
M$10 VGND \$11 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=169000000000P AD=91000000000P PS=1820000U PD=930000U
M$11 X \$11 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=91000000000P AD=108375000000P PS=930000U PD=1010000U
M$12 VGND B1_N \$10 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=108375000000P AD=109200000000P PS=1010000U PD=1360000U
.ENDS sky130_fd_sc_hd__a21bo_2

.SUBCKT sky130_fd_sc_hd__buf_2 VPB A VGND X VPWR VNB
M$1 \$3 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=640000U
+ AS=166400000000P AD=149000000000P PS=1800000U PD=1325000U
M$2 VPWR \$3 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=149000000000P AD=135000000000P PS=1325000U PD=1270000U
M$3 X \$3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=265000000000P PS=1270000U PD=2530000U
M$4 \$3 A VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=109200000000P
+ AD=97000000000P PS=1360000U PD=975000U
M$5 VGND \$3 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=97000000000P
+ AD=87750000000P PS=975000U PD=920000U
M$6 X \$3 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=172250000000P PS=920000U PD=1830000U
.ENDS sky130_fd_sc_hd__buf_2

.SUBCKT sky130_fd_sc_hd__a311o_2 VGND X A3 A2 A1 B1 C1 VPWR VPB VNB
M$1 VPWR \$4 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=135000000000P PS=2520000U PD=1270000U
M$2 X \$4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=240000000000P PS=1270000U PD=1480000U
M$3 VPWR A3 \$13 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=240000000000P AD=170000000000P PS=1480000U PD=1340000U
M$4 \$13 A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=170000000000P AD=185000000000P PS=1340000U PD=1370000U
M$5 VPWR A1 \$13 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=185000000000P AD=210000000000P PS=1370000U PD=1420000U
M$6 \$13 B1 \$15 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=210000000000P AD=210000000000P PS=1420000U PD=1420000U
M$7 \$15 C1 \$4 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=210000000000P AD=260000000000P PS=1420000U PD=2520000U
M$8 VGND \$4 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=169000000000P
+ AD=87750000000P PS=1820000U PD=920000U
M$9 X \$4 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=156000000000P PS=920000U PD=1130000U
M$10 VGND A3 \$6 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=156000000000P AD=110500000000P PS=1130000U PD=990000U
M$11 \$6 A2 \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=110500000000P AD=120250000000P PS=990000U PD=1020000U
M$12 \$5 A1 \$4 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=120250000000P AD=133250000000P PS=1020000U PD=1060000U
M$13 \$4 B1 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=133250000000P AD=139750000000P PS=1060000U PD=1080000U
M$14 VGND C1 \$4 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=139750000000P AD=169000000000P PS=1080000U PD=1820000U
.ENDS sky130_fd_sc_hd__a311o_2

.SUBCKT sky130_fd_sc_hd__and4_2 VPB D C B A VPWR VGND X VNB
M$1 VPWR A \$3 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=109200000000P AD=74550000000P PS=1360000U PD=775000U
M$2 \$3 B VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=74550000000P AD=77700000000P PS=775000U PD=790000U
M$3 VPWR C \$3 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=77700000000P AD=58800000000P PS=790000U PD=700000U
M$4 \$3 D VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=58800000000P AD=279950000000P PS=700000U PD=1615000U
M$5 VPWR \$3 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=279950000000P AD=165000000000P PS=1615000U PD=1330000U
M$6 X \$3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=165000000000P AD=300000000000P PS=1330000U PD=2600000U
M$7 \$3 A \$11 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=109200000000P
+ AD=61950000000P PS=1360000U PD=715000U
M$8 \$11 B \$12 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=61950000000P
+ AD=79800000000P PS=715000U PD=800000U
M$9 \$12 C \$13 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=79800000000P
+ AD=69300000000P PS=800000U PD=750000U
M$10 \$13 D VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=69300000000P AD=175150000000P PS=750000U PD=1265000U
M$11 VGND \$3 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=175150000000P AD=107250000000P PS=1265000U PD=980000U
M$12 X \$3 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=107250000000P AD=195000000000P PS=980000U PD=1900000U
.ENDS sky130_fd_sc_hd__and4_2

.SUBCKT sky130_fd_sc_hd__o221a_2 VGND C1 B1 B2 A2 A1 X VPWR VPB VNB
M$1 \$4 C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=325000000000P AD=165000000000P PS=2650000U PD=1330000U
M$2 VPWR B1 \$13 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=165000000000P AD=112500000000P PS=1330000U PD=1225000U
M$3 \$13 B2 \$4 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=112500000000P AD=387500000000P PS=1225000U PD=1775000U
M$4 \$4 A2 \$14 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=387500000000P AD=105000000000P PS=1775000U PD=1210000U
M$5 \$14 A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=105000000000P AD=165000000000P PS=1210000U PD=1330000U
M$6 VPWR \$4 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=165000000000P AD=135000000000P PS=1330000U PD=1270000U
M$7 X \$4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$8 VGND A2 \$7 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=169000000000P AD=87750000000P PS=1820000U PD=920000U
M$9 \$7 A1 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$10 VGND \$4 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$11 X \$4 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=169000000000P PS=920000U PD=1820000U
M$12 \$4 C1 \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=237250000000P AD=87750000000P PS=2030000U PD=920000U
M$13 \$5 B1 \$7 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$14 \$7 B2 \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=169000000000P PS=920000U PD=1820000U
.ENDS sky130_fd_sc_hd__o221a_2

.SUBCKT sky130_fd_sc_hd__a22oi_2 VGND B2 B1 Y A1 A2 VPWR VPB VNB
M$1 \$10 A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=135000000000P PS=2520000U PD=1270000U
M$2 VPWR A1 \$10 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$3 \$10 A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$4 VPWR A2 \$10 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$5 Y B2 \$10 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=135000000000P PS=2520000U PD=1270000U
M$6 \$10 B2 Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$7 Y B1 \$10 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$8 \$10 B1 Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$9 \$7 A1 Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=169000000000P
+ AD=87750000000P PS=1820000U PD=920000U
M$10 Y A1 \$7 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$11 \$7 A2 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=87750000000P PS=920000U PD=920000U
M$12 VGND A2 \$7 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=169000000000P PS=920000U PD=1820000U
M$13 \$3 B2 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=169000000000P AD=87750000000P PS=1820000U PD=920000U
M$14 VGND B2 \$3 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=87750000000P PS=920000U PD=920000U
M$15 \$3 B1 Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$16 Y B1 \$3 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=169000000000P PS=920000U PD=1820000U
.ENDS sky130_fd_sc_hd__a22oi_2

.SUBCKT sky130_fd_sc_hd__a21o_2 VPB B1 A1 A2 VPWR VGND X VNB
M$1 \$3 B1 \$7 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=265000000000P AD=140000000000P PS=2530000U PD=1280000U
M$2 \$7 A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=157500000000P PS=1280000U PD=1315000U
M$3 VPWR A2 \$7 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=157500000000P AD=260000000000P PS=1315000U PD=2520000U
M$4 VPWR \$3 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=265000000000P AD=140000000000P PS=2530000U PD=1280000U
M$5 X \$3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=265000000000P PS=1280000U PD=2530000U
M$6 VGND \$3 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=172250000000P
+ AD=91000000000P PS=1830000U PD=930000U
M$7 X \$3 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=91000000000P
+ AD=110500000000P PS=930000U PD=990000U
M$8 VGND B1 \$3 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=110500000000P AD=162500000000P PS=990000U PD=1150000U
M$9 \$3 A1 \$11 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=162500000000P AD=123500000000P PS=1150000U PD=1030000U
M$10 \$11 A2 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=123500000000P AD=172250000000P PS=1030000U PD=1830000U
.ENDS sky130_fd_sc_hd__a21o_2

.SUBCKT sky130_fd_sc_hd__o2bb2a_2 VGND X A1_N A2_N B2 B1 VPWR VPB VNB
M$1 VPWR \$4 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=285000000000P AD=135000000000P PS=2570000U PD=1270000U
M$2 X \$4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=154000000000P PS=1270000U PD=1335000U
M$3 VPWR A1_N \$7 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=640000U
+ AS=154000000000P AD=173000000000P PS=1335000U PD=1400000U
M$4 \$7 A2_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=640000U
+ AS=173000000000P AD=227200000000P PS=1400000U PD=1350000U
M$5 VPWR \$7 \$4 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=640000U
+ AS=227200000000P AD=92800000000P PS=1350000U PD=930000U
M$6 \$4 B2 \$13 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=640000U
+ AS=92800000000P AD=86400000000P PS=930000U PD=910000U
M$7 \$13 B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=640000U
+ AS=86400000000P AD=166400000000P PS=910000U PD=1800000U
M$8 \$11 A1_N VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=66150000000P AD=98625000000P PS=735000U PD=980000U
M$9 \$11 A2_N \$7 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=66150000000P AD=109200000000P PS=735000U PD=1360000U
M$10 VGND \$4 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=185250000000P AD=87750000000P PS=1870000U PD=920000U
M$11 X \$4 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=98625000000P PS=920000U PD=980000U
M$12 \$4 \$7 \$8 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=109200000000P AD=56700000000P PS=1360000U PD=690000U
M$13 \$8 B2 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=56700000000P AD=56700000000P PS=690000U PD=690000U
M$14 VGND B1 \$8 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=56700000000P AD=109200000000P PS=690000U PD=1360000U
.ENDS sky130_fd_sc_hd__o2bb2a_2

.SUBCKT sky130_fd_sc_hd__a21oi_2 VPB A1 B1 A2 VPWR Y VGND VNB
M$1 \$7 A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=280000000000P AD=140000000000P PS=2560000U PD=1280000U
M$2 VPWR A1 \$7 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$3 \$7 A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=135000000000P PS=1280000U PD=1270000U
M$4 VPWR A2 \$7 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$5 \$7 B1 Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$6 Y B1 \$7 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=360000000000P PS=1270000U PD=2720000U
M$7 VGND A2 \$10 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=185250000000P AD=89375000000P PS=1870000U PD=925000U
M$8 \$10 A1 Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=89375000000P
+ AD=91000000000P PS=925000U PD=930000U
M$9 Y A1 \$11 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=91000000000P
+ AD=68250000000P PS=930000U PD=860000U
M$10 \$11 A2 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=68250000000P AD=107250000000P PS=860000U PD=980000U
M$11 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=107250000000P
+ AD=87750000000P PS=980000U PD=920000U
M$12 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=260000000000P PS=920000U PD=2100000U
.ENDS sky130_fd_sc_hd__a21oi_2

.SUBCKT sky130_fd_sc_hd__a2bb2o_2 VGND X B1 A1_N A2_N B2 VPWR VPB VNB
M$1 \$7 \$4 \$12 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=640000U
+ AS=166400000000P AD=97600000000P PS=1800000U PD=945000U
M$2 \$12 B2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=640000U
+ AS=97600000000P AD=86400000000P PS=945000U PD=910000U
M$3 VPWR B1 \$12 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=640000U
+ AS=86400000000P AD=166400000000P PS=910000U PD=1800000U
M$4 \$13 A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=640000U
+ AS=67200000000P AD=186000000000P PS=850000U PD=1435000U
M$5 \$13 A2_N \$4 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=640000U
+ AS=67200000000P AD=169600000000P PS=850000U PD=1810000U
M$6 VPWR \$7 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=265000000000P AD=135000000000P PS=2530000U PD=1270000U
M$7 X \$7 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=186000000000P PS=1270000U PD=1435000U
M$8 \$4 A1_N VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=56700000000P AD=120100000000P PS=690000U PD=1085000U
M$9 \$4 A2_N VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=56700000000P AD=141750000000P PS=690000U PD=1095000U
M$10 VGND \$4 \$7 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=141750000000P AD=56700000000P PS=1095000U PD=690000U
M$11 \$7 B2 \$6 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=56700000000P
+ AD=56700000000P PS=690000U PD=690000U
M$12 \$6 B1 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=56700000000P AD=109200000000P PS=690000U PD=1360000U
M$13 VGND \$7 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=172250000000P AD=87750000000P PS=1830000U PD=920000U
M$14 X \$7 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=120100000000P PS=920000U PD=1085000U
.ENDS sky130_fd_sc_hd__a2bb2o_2

.SUBCKT sky130_fd_sc_hd__o21a_2 VPB B1 A2 A1 VGND VPWR X VNB
M$1 VPWR \$3 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=137500000000P PS=2520000U PD=1275000U
M$2 X \$3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=137500000000P AD=400000000000P PS=1275000U PD=1800000U
M$3 VPWR B1 \$3 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=400000000000P AD=140000000000P PS=1800000U PD=1280000U
M$4 \$3 A2 \$11 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=160000000000P PS=1280000U PD=1320000U
M$5 \$11 A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=160000000000P AD=265000000000P PS=1320000U PD=2530000U
M$6 VGND \$3 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=169000000000P
+ AD=89375000000P PS=1820000U PD=925000U
M$7 X \$3 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=89375000000P
+ AD=172250000000P PS=925000U PD=1830000U
M$8 \$3 B1 \$10 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=172250000000P AD=91000000000P PS=1830000U PD=930000U
M$9 \$10 A2 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=91000000000P AD=104000000000P PS=930000U PD=970000U
M$10 VGND A1 \$10 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=104000000000P AD=172250000000P PS=970000U PD=1830000U
.ENDS sky130_fd_sc_hd__o21a_2

.SUBCKT sky130_fd_sc_hd__and3_2 VPB A B C VGND VPWR X VNB
M$1 \$6 C VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=74375000000P AD=150750000000P PS=815000U PD=1345000U
M$2 \$6 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=109200000000P AD=56700000000P PS=1360000U PD=690000U
M$3 VPWR B \$6 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=56700000000P AD=74375000000P PS=690000U PD=815000U
M$4 VPWR \$6 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=150750000000P AD=135000000000P PS=1345000U PD=1270000U
M$5 X \$6 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$6 \$6 A \$11 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=109200000000P
+ AD=44100000000P PS=1360000U PD=630000U
M$7 \$11 B \$10 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=44100000000P
+ AD=53550000000P PS=630000U PD=675000U
M$8 \$10 C VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=53550000000P
+ AD=130400000000P PS=675000U PD=1105000U
M$9 VGND \$6 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=130400000000P
+ AD=87750000000P PS=1105000U PD=920000U
M$10 X \$6 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=178750000000P PS=920000U PD=1850000U
.ENDS sky130_fd_sc_hd__and3_2

.SUBCKT sky130_fd_sc_hd__or4_2 VPB D C B A VGND VPWR X VNB
M$1 \$7 D \$11 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=109200000000P AD=69300000000P PS=1360000U PD=750000U
M$2 \$11 C \$12 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=69300000000P AD=44100000000P PS=750000U PD=630000U
M$3 \$12 B \$13 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=44100000000P AD=69300000000P PS=630000U PD=750000U
M$4 \$13 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=69300000000P AD=148250000000P PS=750000U PD=1340000U
M$5 VPWR \$7 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=148250000000P AD=135000000000P PS=1340000U PD=1270000U
M$6 X \$7 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=305000000000P PS=1270000U PD=2610000U
M$7 VGND D \$7 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=109200000000P
+ AD=69300000000P PS=1360000U PD=750000U
M$8 \$7 C VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=69300000000P
+ AD=56700000000P PS=750000U PD=690000U
M$9 VGND B \$7 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=56700000000P
+ AD=56700000000P PS=690000U PD=690000U
M$10 \$7 A VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=56700000000P
+ AD=101875000000P PS=690000U PD=990000U
M$11 VGND \$7 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=101875000000P AD=87750000000P PS=990000U PD=920000U
M$12 X \$7 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=198250000000P PS=920000U PD=1910000U
.ENDS sky130_fd_sc_hd__or4_2

.SUBCKT sky130_fd_sc_hd__conb_1 VPB HI|VPWR LO|VGND VNB
R$1 LO|VGND LO|VGND 0
R$2 HI|VPWR HI|VPWR 0
.ENDS sky130_fd_sc_hd__conb_1

.SUBCKT sky130_fd_sc_hd__clkinv_2 VPB A Y VPWR VGND VNB
M$1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=265000000000P AD=140000000000P PS=2530000U PD=1280000U
M$2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$3 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=265000000000P PS=1280000U PD=2530000U
M$4 VGND A Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=111300000000P
+ AD=58800000000P PS=1370000U PD=700000U
M$5 Y A VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=109200000000P PS=700000U PD=1360000U
.ENDS sky130_fd_sc_hd__clkinv_2

.SUBCKT sky130_fd_sc_hd__clkinv_8 VGND Y A VPWR VPB VNB
M$1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=135000000000P PS=2520000U PD=1270000U
M$2 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=137500000000P PS=1270000U PD=1275000U
M$3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=137500000000P AD=135000000000P PS=1275000U PD=1270000U
M$4 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$5 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$6 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$7 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$9 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$10 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$11 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$12 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$13 VGND A Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=111300000000P
+ AD=58800000000P PS=1370000U PD=700000U
M$14 Y A VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=58800000000P PS=700000U PD=700000U
M$15 VGND A Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=58800000000P PS=700000U PD=700000U
M$16 Y A VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=58800000000P PS=700000U PD=700000U
M$17 VGND A Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=58800000000P PS=700000U PD=700000U
M$18 Y A VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=58800000000P PS=700000U PD=700000U
M$19 VGND A Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=58800000000P PS=700000U PD=700000U
M$20 Y A VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=111300000000P PS=700000U PD=1370000U
.ENDS sky130_fd_sc_hd__clkinv_8

.SUBCKT sky130_fd_sc_hd__einvp_1 VPB A TE VPWR Z VGND VNB
M$1 \$8 TE VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=109200000000P AD=320750000000P PS=1360000U PD=1685000U
M$2 VPWR \$8 \$9 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=320750000000P AD=182500000000P PS=1685000U PD=1365000U
M$3 \$9 A Z VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=182500000000P AD=270000000000P PS=1365000U PD=2540000U
M$4 \$8 TE VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=109200000000P AD=97000000000P PS=1360000U PD=975000U
M$5 VGND TE \$10 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=97000000000P AD=235625000000P PS=975000U PD=1375000U
M$6 \$10 A Z VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=235625000000P
+ AD=175500000000P PS=1375000U PD=1840000U
.ENDS sky130_fd_sc_hd__einvp_1

.SUBCKT sky130_fd_sc_hd__nand2_2 VPB A B VPWR Y VGND VNB
M$1 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=135000000000P PS=2520000U PD=1270000U
M$2 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$4 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$5 \$6 B VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=169000000000P
+ AD=87750000000P PS=1820000U PD=920000U
M$6 VGND B \$6 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$7 \$6 A Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$8 Y A \$6 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=169000000000P PS=920000U PD=1820000U
.ENDS sky130_fd_sc_hd__nand2_2

.SUBCKT sky130_fd_sc_hd__and2_2 VPB A B VPWR X VGND VNB
M$1 VPWR A \$5 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=117600000000P AD=56700000000P PS=1400000U PD=690000U
M$2 \$5 B VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=56700000000P AD=166550000000P PS=690000U PD=1390000U
M$3 VPWR \$5 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=166550000000P AD=195000000000P PS=1390000U PD=1390000U
M$4 X \$5 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=195000000000P AD=380000000000P PS=1390000U PD=2760000U
M$5 \$5 A \$9 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=117600000000P
+ AD=56700000000P PS=1400000U PD=690000U
M$6 \$9 B VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=56700000000P
+ AD=111800000000P PS=690000U PD=1040000U
M$7 VGND \$5 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=111800000000P
+ AD=126750000000P PS=1040000U PD=1040000U
M$8 X \$5 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=126750000000P
+ AD=247000000000P PS=1040000U PD=2060000U
.ENDS sky130_fd_sc_hd__and2_2

.SUBCKT sky130_fd_sc_hd__a32o_2 VGND X B2 A2 B1 A1 A3 VPWR VPB VNB
M$1 \$14 B2 \$5 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=135000000000P PS=2520000U PD=1270000U
M$2 \$5 B1 \$14 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$3 \$14 A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=215000000000P PS=1270000U PD=1430000U
M$4 VPWR A2 \$14 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=215000000000P AD=135000000000P PS=1430000U PD=1270000U
M$5 \$14 A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$6 X \$5 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=135000000000P PS=2520000U PD=1270000U
M$7 VPWR \$5 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$8 VGND \$5 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=169000000000P
+ AD=87750000000P PS=1820000U PD=920000U
M$9 X \$5 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=209625000000P PS=920000U PD=1295000U
M$10 VGND B2 \$11 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=209625000000P AD=115375000000P PS=1295000U PD=1005000U
M$11 \$11 B1 \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=115375000000P AD=107250000000P PS=1005000U PD=980000U
M$12 \$5 A1 \$12 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=107250000000P AD=139750000000P PS=980000U PD=1080000U
M$13 \$12 A2 \$10 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=139750000000P AD=87750000000P PS=1080000U PD=920000U
M$14 \$10 A3 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=169000000000P PS=920000U PD=1820000U
.ENDS sky130_fd_sc_hd__a32o_2

.SUBCKT sky130_fd_sc_hd__a31o_2 VPB B1 A1 A2 A3 X VPWR VGND VNB
M$1 VPWR \$11 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=135000000000P PS=2520000U PD=1270000U
M$2 X \$11 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$3 VPWR A3 \$10 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$4 \$10 A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=165000000000P PS=1270000U PD=1330000U
M$5 VPWR A1 \$10 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=165000000000P AD=165000000000P PS=1330000U PD=1330000U
M$6 \$10 B1 \$11 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=165000000000P AD=320000000000P PS=1330000U PD=2640000U
M$7 VGND \$11 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=169000000000P AD=87750000000P PS=1820000U PD=920000U
M$8 X \$11 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$9 VGND A3 \$12 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=87750000000P PS=920000U PD=920000U
M$10 \$12 A2 \$13 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=107250000000P PS=920000U PD=980000U
M$11 \$13 A1 \$11 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=107250000000P AD=126750000000P PS=980000U PD=1040000U
M$12 \$11 B1 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=126750000000P AD=169000000000P PS=1040000U PD=1820000U
.ENDS sky130_fd_sc_hd__a31o_2

.SUBCKT sky130_fd_sc_hd__o32a_2 VGND X A1 A2 A3 B2 B1 VPWR VPB VNB
M$1 VPWR \$5 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=135000000000P PS=2520000U PD=1270000U
M$2 X \$5 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=305000000000P PS=1270000U PD=1610000U
M$3 VPWR A1 \$13 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=305000000000P AD=135000000000P PS=1610000U PD=1270000U
M$4 \$13 A2 \$12 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=215000000000P PS=1270000U PD=1430000U
M$5 \$12 A3 \$5 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=215000000000P AD=135000000000P PS=1430000U PD=1270000U
M$6 \$5 B2 \$14 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=190000000000P PS=1270000U PD=1380000U
M$7 \$14 B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=190000000000P AD=330000000000P PS=1380000U PD=2660000U
M$8 VGND \$5 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=169000000000P
+ AD=87750000000P PS=1820000U PD=920000U
M$9 X \$5 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=198250000000P PS=920000U PD=1260000U
M$10 VGND A1 \$4 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=198250000000P AD=87750000000P PS=1260000U PD=920000U
M$11 \$4 A2 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=139750000000P PS=920000U PD=1080000U
M$12 VGND A3 \$4 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=139750000000P AD=87750000000P PS=1080000U PD=920000U
M$13 \$4 B2 \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=123500000000P PS=920000U PD=1030000U
M$14 \$5 B1 \$4 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=123500000000P AD=214500000000P PS=1030000U PD=1960000U
.ENDS sky130_fd_sc_hd__o32a_2

.SUBCKT sky130_fd_sc_hd__o31a_2 VPB A1 A2 A3 B1 VPWR VGND X VNB
M$1 VPWR \$11 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=405000000000P AD=175000000000P PS=2810000U PD=1350000U
M$2 X \$11 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=175000000000P AD=195000000000P PS=1350000U PD=1390000U
M$3 VPWR A1 \$13 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=195000000000P AD=135000000000P PS=1390000U PD=1270000U
M$4 \$13 A2 \$12 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=165000000000P PS=1270000U PD=1330000U
M$5 \$12 A3 \$11 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=165000000000P AD=212500000000P PS=1330000U PD=1425000U
M$6 \$11 B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=212500000000P AD=340000000000P PS=1425000U PD=2680000U
M$7 VGND \$11 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=263250000000P AD=113750000000P PS=2110000U PD=1000000U
M$8 X \$11 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=113750000000P AD=126750000000P PS=1000000U PD=1040000U
M$9 VGND A1 \$10 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=126750000000P AD=87750000000P PS=1040000U PD=920000U
M$10 \$10 A2 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=107250000000P PS=920000U PD=980000U
M$11 VGND A3 \$10 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=107250000000P AD=107250000000P PS=980000U PD=980000U
M$12 \$10 B1 \$11 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=107250000000P AD=201500000000P PS=980000U PD=1920000U
.ENDS sky130_fd_sc_hd__o31a_2

.SUBCKT sky130_fd_sc_hd__nor2_2 VPB A B VGND VPWR Y VNB
M$1 \$6 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=280000000000P AD=135000000000P PS=2560000U PD=1270000U
M$2 VPWR A \$6 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$3 \$6 B Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$4 Y B \$6 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$5 VGND A Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=182000000000P
+ AD=87750000000P PS=1860000U PD=920000U
M$6 Y A VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$7 VGND B Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$8 Y B VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=169000000000P PS=920000U PD=1820000U
.ENDS sky130_fd_sc_hd__nor2_2

.SUBCKT sky130_fd_sc_hd__decap_8 VPB VGND VPWR VNB
M$1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=2890000U W=870000U
+ AS=226200000000P AD=226200000000P PS=2260000U PD=2260000U
M$2 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 L=2890000U W=550000U
+ AS=143000000000P AD=143000000000P PS=1620000U PD=1620000U
.ENDS sky130_fd_sc_hd__decap_8

.SUBCKT sky130_fd_sc_hd__clkinv_1 VPB A VPWR VGND Y VNB
M$1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=840000U
+ AS=218400000000P AD=113400000000P PS=2200000U PD=1110000U
M$2 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=840000U
+ AS=113400000000P AD=235200000000P PS=1110000U PD=2240000U
M$3 Y A VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=109200000000P
+ AD=119700000000P PS=1360000U PD=1410000U
.ENDS sky130_fd_sc_hd__clkinv_1

.SUBCKT sky130_fd_sc_hd__decap_12 VPB VGND VPWR VNB
M$1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=4730000U W=870000U
+ AS=226200000000P AD=226200000000P PS=2260000U PD=2260000U
M$2 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 L=4730000U W=550000U
+ AS=143000000000P AD=143000000000P PS=1620000U PD=1620000U
.ENDS sky130_fd_sc_hd__decap_12

.SUBCKT sky130_fd_sc_hd__einvn_8 VGND A TE_B Z VPWR VPB VNB
M$1 \$6 TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=160250000000P PS=2520000U PD=1325000U
M$2 VPWR TE_B \$8 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=940000U
+ AS=160250000000P AD=126900000000P PS=1325000U PD=1210000U
M$3 \$8 TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=940000U
+ AS=126900000000P AD=126900000000P PS=1210000U PD=1210000U
M$4 VPWR TE_B \$8 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=940000U
+ AS=126900000000P AD=126900000000P PS=1210000U PD=1210000U
M$5 \$8 TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=940000U
+ AS=126900000000P AD=126900000000P PS=1210000U PD=1210000U
M$6 VPWR TE_B \$8 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=940000U
+ AS=126900000000P AD=126900000000P PS=1210000U PD=1210000U
M$7 \$8 TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=940000U
+ AS=126900000000P AD=126900000000P PS=1210000U PD=1210000U
M$8 VPWR TE_B \$8 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=940000U
+ AS=126900000000P AD=126900000000P PS=1210000U PD=1210000U
M$9 \$8 TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=940000U
+ AS=126900000000P AD=244400000000P PS=1210000U PD=2400000U
M$10 \$8 A Z VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=135000000000P PS=2520000U PD=1270000U
M$11 Z A \$8 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$12 \$8 A Z VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$13 Z A \$8 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$14 \$8 A Z VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$15 Z A \$8 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$16 \$8 A Z VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$17 Z A \$8 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$18 \$5 \$6 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=169000000000P AD=87750000000P PS=1820000U PD=920000U
M$19 VGND \$6 \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=87750000000P PS=920000U PD=920000U
M$20 \$5 \$6 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=87750000000P PS=920000U PD=920000U
M$21 VGND \$6 \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=87750000000P PS=920000U PD=920000U
M$22 \$5 \$6 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=87750000000P PS=920000U PD=920000U
M$23 VGND \$6 \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=87750000000P PS=920000U PD=920000U
M$24 \$5 \$6 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=87750000000P PS=920000U PD=920000U
M$25 VGND \$6 \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=105625000000P PS=920000U PD=975000U
M$26 \$5 A Z VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=105625000000P
+ AD=87750000000P PS=975000U PD=920000U
M$27 Z A \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$28 \$5 A Z VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$29 Z A \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$30 \$5 A Z VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$31 Z A \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$32 \$5 A Z VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$33 Z A \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=182000000000P PS=920000U PD=1860000U
M$34 \$6 TE_B VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=169000000000P AD=169000000000P PS=1820000U PD=1820000U
.ENDS sky130_fd_sc_hd__einvn_8

.SUBCKT sky130_fd_sc_hd__clkbuf_2 VPB A VPWR VGND X VNB
M$1 \$6 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=265000000000P AD=162500000000P PS=2530000U PD=1325000U
M$2 VPWR \$6 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=162500000000P AD=135000000000P PS=1325000U PD=1270000U
M$3 X \$6 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$4 \$6 A VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=111300000000P
+ AD=68250000000P PS=1370000U PD=745000U
M$5 VGND \$6 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=68250000000P
+ AD=56700000000P PS=745000U PD=690000U
M$6 X \$6 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=56700000000P
+ AD=109200000000P PS=690000U PD=1360000U
.ENDS sky130_fd_sc_hd__clkbuf_2

.SUBCKT sky130_fd_sc_hd__or3_2 VPB B A C VPWR VGND X VNB
M$1 \$9 C \$11 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=109200000000P AD=44100000000P PS=1360000U PD=630000U
M$2 \$11 B \$10 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=44100000000P AD=69300000000P PS=630000U PD=750000U
M$3 \$10 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=69300000000P AD=148250000000P PS=750000U PD=1340000U
M$4 VPWR \$9 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=148250000000P AD=135000000000P PS=1340000U PD=1270000U
M$5 X \$9 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=315000000000P PS=1270000U PD=2630000U
M$6 \$9 C VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=109200000000P
+ AD=56700000000P PS=1360000U PD=690000U
M$7 VGND B \$9 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=56700000000P
+ AD=56700000000P PS=690000U PD=690000U
M$8 \$9 A VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=56700000000P
+ AD=101875000000P PS=690000U PD=990000U
M$9 VGND \$9 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=101875000000P
+ AD=87750000000P PS=990000U PD=920000U
M$10 X \$9 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=185250000000P PS=920000U PD=1870000U
.ENDS sky130_fd_sc_hd__or3_2

.SUBCKT sky130_fd_sc_hd__a221o_2 VGND C1 B2 B1 A1 A2 X VPWR VPB VNB
M$1 VPWR A1 \$14 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=165000000000P PS=2520000U PD=1330000U
M$2 \$14 A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=165000000000P AD=157500000000P PS=1330000U PD=1315000U
M$3 VPWR \$3 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=157500000000P AD=135000000000P PS=1315000U PD=1270000U
M$4 X \$3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=285000000000P PS=1270000U PD=2570000U
M$5 \$3 C1 \$13 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=135000000000P PS=2520000U PD=1270000U
M$6 \$13 B2 \$14 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$7 \$14 B1 \$13 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$8 \$3 A1 \$11 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=169000000000P AD=107250000000P PS=1820000U PD=980000U
M$9 \$11 A2 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=107250000000P AD=102375000000P PS=980000U PD=965000U
M$10 VGND \$3 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=102375000000P AD=87750000000P PS=965000U PD=920000U
M$11 X \$3 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=185250000000P PS=920000U PD=1870000U
M$12 \$3 C1 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=169000000000P AD=107250000000P PS=1820000U PD=980000U
M$13 VGND B2 \$10 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=107250000000P AD=68250000000P PS=980000U PD=860000U
M$14 \$10 B1 \$3 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=68250000000P AD=169000000000P PS=860000U PD=1820000U
.ENDS sky130_fd_sc_hd__a221o_2

.SUBCKT sky130_fd_sc_hd__clkbuf_1 VPB A X VGND VPWR VNB
M$1 X \$3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=790000U
+ AS=205400000000P AD=114550000000P PS=2100000U PD=1080000U
M$2 VPWR A \$3 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=790000U
+ AS=114550000000P AD=205400000000P PS=1080000U PD=2100000U
M$3 X \$3 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=520000U AS=135200000000P
+ AD=75400000000P PS=1560000U PD=810000U
M$4 VGND A \$3 VNB sky130_fd_pr__nfet_01v8 L=150000U W=520000U AS=75400000000P
+ AD=135200000000P PS=810000U PD=1560000U
.ENDS sky130_fd_sc_hd__clkbuf_1

.SUBCKT sky130_fd_sc_hd__einvp_2 VPB TE A Z VPWR VGND VNB
M$1 \$8 TE VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=640000U
+ AS=166400000000P AD=166400000000P PS=1800000U PD=1800000U
M$2 \$5 \$8 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=940000U
+ AS=244400000000P AD=126900000000P PS=2400000U PD=1210000U
M$3 VPWR \$8 \$5 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=940000U
+ AS=126900000000P AD=160250000000P PS=1210000U PD=1325000U
M$4 \$5 A Z VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=160250000000P AD=135000000000P PS=1325000U PD=1270000U
M$5 Z A \$5 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$6 \$8 TE VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=109200000000P AD=97000000000P PS=1360000U PD=975000U
M$7 VGND TE \$7 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=97000000000P
+ AD=87750000000P PS=975000U PD=920000U
M$8 \$7 TE VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=169000000000P PS=920000U PD=1820000U
M$9 \$7 A Z VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=169000000000P
+ AD=87750000000P PS=1820000U PD=920000U
M$10 Z A \$7 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=169000000000P PS=920000U PD=1820000U
.ENDS sky130_fd_sc_hd__einvp_2

.SUBCKT sky130_fd_sc_hd__o311a_2 VGND X A1 A2 A3 B1 C1 VPWR VPB VNB
M$1 VPWR \$5 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=320000000000P AD=135000000000P PS=2640000U PD=1270000U
M$2 X \$5 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=312500000000P PS=1270000U PD=1625000U
M$3 VPWR A1 \$15 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=312500000000P AD=175000000000P PS=1625000U PD=1350000U
M$4 \$15 A2 \$14 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=175000000000P AD=210000000000P PS=1350000U PD=1420000U
M$5 \$14 A3 \$5 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=210000000000P AD=137500000000P PS=1420000U PD=1275000U
M$6 \$5 B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=137500000000P AD=150000000000P PS=1275000U PD=1300000U
M$7 VPWR C1 \$5 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=150000000000P AD=260000000000P PS=1300000U PD=2520000U
M$8 VGND \$5 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=208000000000P
+ AD=87750000000P PS=1940000U PD=920000U
M$9 X \$5 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=203125000000P PS=920000U PD=1275000U
M$10 VGND A1 \$4 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=203125000000P AD=113750000000P PS=1275000U PD=1000000U
M$11 \$4 A2 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=113750000000P AD=136500000000P PS=1000000U PD=1070000U
M$12 VGND A3 \$4 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=136500000000P AD=118625000000P PS=1070000U PD=1015000U
M$13 \$4 B1 \$11 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=118625000000P AD=68250000000P PS=1015000U PD=860000U
M$14 \$11 C1 \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=68250000000P AD=169000000000P PS=860000U PD=1820000U
.ENDS sky130_fd_sc_hd__o311a_2

.SUBCKT sky130_fd_sc_hd__o21ai_2 VPB A1 A2 B1 VGND Y VPWR VNB
M$1 VPWR A1 \$7 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=265000000000P AD=140000000000P PS=2530000U PD=1280000U
M$2 \$7 A2 Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$3 Y A2 \$7 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=175000000000P PS=1280000U PD=1350000U
M$4 \$7 A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=175000000000P AD=160000000000P PS=1350000U PD=1320000U
M$5 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=160000000000P AD=140000000000P PS=1320000U PD=1280000U
M$6 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=265000000000P PS=1280000U PD=2530000U
M$7 \$6 A1 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=172250000000P AD=91000000000P PS=1830000U PD=930000U
M$8 VGND A2 \$6 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=91000000000P
+ AD=91000000000P PS=930000U PD=930000U
M$9 \$6 A2 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=91000000000P
+ AD=126750000000P PS=930000U PD=1040000U
M$10 VGND A1 \$6 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=126750000000P AD=91000000000P PS=1040000U PD=930000U
M$11 \$6 B1 Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=91000000000P
+ AD=91000000000P PS=930000U PD=930000U
M$12 Y B1 \$6 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=91000000000P
+ AD=172250000000P PS=930000U PD=1830000U
.ENDS sky130_fd_sc_hd__o21ai_2

.SUBCKT sky130_fd_sc_hd__o22a_2 VPB B1 B2 A2 A1 VPWR X VGND VNB
M$1 VPWR \$3 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=280000000000P AD=135000000000P PS=2560000U PD=1270000U
M$2 X \$3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=390000000000P PS=1270000U PD=1780000U
M$3 VPWR B1 \$12 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=390000000000P AD=105000000000P PS=1780000U PD=1210000U
M$4 \$12 B2 \$3 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=105000000000P AD=235000000000P PS=1210000U PD=1470000U
M$5 \$3 A2 \$13 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=235000000000P AD=105000000000P PS=1470000U PD=1210000U
M$6 \$13 A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=105000000000P AD=280000000000P PS=1210000U PD=2560000U
M$7 VGND \$3 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=169000000000P
+ AD=87750000000P PS=1820000U PD=920000U
M$8 X \$3 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=169000000000P PS=920000U PD=1820000U
M$9 \$10 B1 \$3 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=169000000000P AD=87750000000P PS=1820000U PD=920000U
M$10 \$3 B2 \$10 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=123500000000P PS=920000U PD=1030000U
M$11 \$10 A2 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=123500000000P AD=87750000000P PS=1030000U PD=920000U
M$12 VGND A1 \$10 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=169000000000P PS=920000U PD=1820000U
.ENDS sky130_fd_sc_hd__o22a_2

.SUBCKT sky130_fd_sc_hd__or2_2 VPB A B X VPWR VGND VNB
M$1 \$4 B \$9 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=109200000000P AD=44100000000P PS=1360000U PD=630000U
M$2 \$9 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=44100000000P AD=155750000000P PS=630000U PD=1355000U
M$3 VPWR \$4 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=155750000000P AD=135000000000P PS=1355000U PD=1270000U
M$4 X \$4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$5 VGND B \$4 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=109200000000P
+ AD=56700000000P PS=1360000U PD=690000U
M$6 \$4 A VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=56700000000P
+ AD=106750000000P PS=690000U PD=1005000U
M$7 VGND \$4 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=106750000000P
+ AD=87750000000P PS=1005000U PD=920000U
M$8 X \$4 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=169000000000P PS=920000U PD=1820000U
.ENDS sky130_fd_sc_hd__or2_2

.SUBCKT sky130_fd_sc_hd__decap_4 VPB VGND VPWR VNB
M$1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=1050000U W=870000U
+ AS=226200000000P AD=226200000000P PS=2260000U PD=2260000U
M$2 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 L=1050000U W=550000U
+ AS=143000000000P AD=143000000000P PS=1620000U PD=1620000U
.ENDS sky130_fd_sc_hd__decap_4

.SUBCKT sky130_fd_sc_hd__buf_1 VPB A X VGND VPWR VNB
M$1 \$3 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=790000U
+ AS=205400000000P AD=114550000000P PS=2100000U PD=1080000U
M$2 VPWR \$3 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=790000U
+ AS=114550000000P AD=205400000000P PS=1080000U PD=2100000U
M$3 \$3 A VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=520000U AS=135200000000P
+ AD=75400000000P PS=1560000U PD=810000U
M$4 VGND \$3 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=520000U AS=75400000000P
+ AD=135200000000P PS=810000U PD=1560000U
.ENDS sky130_fd_sc_hd__buf_1

.SUBCKT sky130_fd_sc_hd__o41a_2 VGND X B1 A4 A3 A2 A1 VPWR VPB VNB
M$1 VPWR \$4 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=135000000000P PS=2520000U PD=1270000U
M$2 X \$4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=305000000000P PS=1270000U PD=1610000U
M$3 VPWR B1 \$4 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=305000000000P AD=302500000000P PS=1610000U PD=1605000U
M$4 \$4 A4 \$13 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=302500000000P AD=177500000000P PS=1605000U PD=1355000U
M$5 \$13 A3 \$14 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=177500000000P AD=175000000000P PS=1355000U PD=1350000U
M$6 \$14 A2 \$15 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=175000000000P AD=175000000000P PS=1350000U PD=1350000U
M$7 \$15 A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=175000000000P AD=410000000000P PS=1350000U PD=2820000U
M$8 VGND \$4 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=169000000000P
+ AD=87750000000P PS=1820000U PD=920000U
M$9 X \$4 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=169000000000P PS=920000U PD=1820000U
M$10 \$4 B1 \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=208000000000P AD=118625000000P PS=1940000U PD=1015000U
M$11 \$5 A4 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=118625000000P AD=115375000000P PS=1015000U PD=1005000U
M$12 VGND A3 \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=115375000000P AD=113750000000P PS=1005000U PD=1000000U
M$13 \$5 A2 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=113750000000P AD=113750000000P PS=1000000U PD=1000000U
M$14 VGND A1 \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=113750000000P AD=266500000000P PS=1000000U PD=2120000U
.ENDS sky130_fd_sc_hd__o41a_2

.SUBCKT sky130_fd_sc_hd__einvn_4 VGND A Z TE_B VPWR VPB VNB
M$1 \$8 A Z VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=135000000000P PS=2520000U PD=1270000U
M$2 Z A \$8 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$3 \$8 A Z VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$4 Z A \$8 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$5 \$4 TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=160250000000P PS=2520000U PD=1325000U
M$6 VPWR TE_B \$8 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=940000U
+ AS=160250000000P AD=126900000000P PS=1325000U PD=1210000U
M$7 \$8 TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=940000U
+ AS=126900000000P AD=126900000000P PS=1210000U PD=1210000U
M$8 VPWR TE_B \$8 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=940000U
+ AS=126900000000P AD=126900000000P PS=1210000U PD=1210000U
M$9 \$8 TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=940000U
+ AS=126900000000P AD=244400000000P PS=1210000U PD=2400000U
M$10 \$5 \$4 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=169000000000P AD=87750000000P PS=1820000U PD=920000U
M$11 VGND \$4 \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=87750000000P PS=920000U PD=920000U
M$12 \$5 \$4 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=87750000000P PS=920000U PD=920000U
M$13 VGND \$4 \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=105625000000P PS=920000U PD=975000U
M$14 \$5 A Z VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=105625000000P
+ AD=87750000000P PS=975000U PD=920000U
M$15 Z A \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$16 \$5 A Z VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$17 Z A \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=182000000000P PS=920000U PD=1860000U
M$18 \$4 TE_B VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=169000000000P AD=169000000000P PS=1820000U PD=1820000U
.ENDS sky130_fd_sc_hd__einvn_4

.SUBCKT sky130_fd_sc_hd__mux2_1 VPB S A1 A0 X VPWR VGND VNB
M$1 \$11 S VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=76650000000P AD=158350000000P PS=785000U PD=1395000U
M$2 \$11 A0 \$8 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=76650000000P AD=193200000000P PS=785000U PD=1340000U
M$3 \$8 A1 \$12 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=193200000000P AD=44100000000P PS=1340000U PD=630000U
M$4 \$12 \$4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=44100000000P AD=69300000000P PS=630000U PD=750000U
M$5 VPWR S \$4 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=69300000000P AD=117600000000P PS=750000U PD=1400000U
M$6 X \$8 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=158350000000P PS=2520000U PD=1395000U
M$7 \$13 S VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=69300000000P
+ AD=112850000000P PS=750000U PD=1045000U
M$8 \$13 A1 \$8 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=69300000000P
+ AD=99750000000P PS=750000U PD=895000U
M$9 \$8 A0 \$14 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=99750000000P
+ AD=69300000000P PS=895000U PD=750000U
M$10 \$14 \$4 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=69300000000P AD=144900000000P PS=750000U PD=1110000U
M$11 VGND S \$4 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=144900000000P AD=109200000000P PS=1110000U PD=1360000U
M$12 X \$8 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=169000000000P AD=112850000000P PS=1820000U PD=1045000U
.ENDS sky130_fd_sc_hd__mux2_1

.SUBCKT sky130_fd_sc_hd__decap_3 VPB VGND VPWR VNB
M$1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=590000U W=870000U
+ AS=226200000000P AD=226200000000P PS=2260000U PD=2260000U
M$2 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 L=590000U W=550000U
+ AS=143000000000P AD=143000000000P PS=1620000U PD=1620000U
.ENDS sky130_fd_sc_hd__decap_3

.SUBCKT sky130_fd_sc_hd__o211a_2 VPB C1 B1 A2 A1 VPWR VGND X VNB
M$1 \$7 C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=265000000000P AD=140000000000P PS=2530000U PD=1280000U
M$2 VPWR B1 \$7 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=367500000000P PS=1280000U PD=1735000U
M$3 \$7 A2 \$12 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=367500000000P AD=105000000000P PS=1735000U PD=1210000U
M$4 \$12 A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=105000000000P AD=195000000000P PS=1210000U PD=1390000U
M$5 VPWR \$7 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=195000000000P AD=140000000000P PS=1390000U PD=1280000U
M$6 X \$7 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=265000000000P PS=1280000U PD=2530000U
M$7 VGND A2 \$9 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=165350000000P AD=91000000000P PS=1820000U PD=930000U
M$8 \$9 A1 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=91000000000P
+ AD=104000000000P PS=930000U PD=970000U
M$9 VGND \$7 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=104000000000P
+ AD=91000000000P PS=970000U PD=930000U
M$10 X \$7 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=91000000000P
+ AD=230750000000P PS=930000U PD=2010000U
M$11 \$7 C1 \$13 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=172250000000P AD=68250000000P PS=1830000U PD=860000U
M$12 \$13 B1 \$9 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=68250000000P AD=165350000000P PS=860000U PD=1820000U
.ENDS sky130_fd_sc_hd__o211a_2

.SUBCKT sky130_fd_sc_hd__inv_2 VPB A VGND VPWR Y VNB
M$1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=135000000000P PS=2520000U PD=1270000U
M$2 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$3 VGND A Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=169000000000P
+ AD=87750000000P PS=1820000U PD=920000U
M$4 Y A VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=169000000000P PS=920000U PD=1820000U
.ENDS sky130_fd_sc_hd__inv_2

.SUBCKT sky130_fd_sc_hd__decap_6 VPB VPWR VGND VNB
M$1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=1970000U W=870000U
+ AS=226200000000P AD=226200000000P PS=2260000U PD=2260000U
M$2 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 L=1970000U W=550000U
+ AS=143000000000P AD=143000000000P PS=1620000U PD=1620000U
.ENDS sky130_fd_sc_hd__decap_6

.SUBCKT sky130_fd_sc_hd__o221ai_2 VGND C1 Y B1 B2 A1 A2 VPWR VPB VNB
M$1 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=135000000000P PS=2520000U PD=1270000U
M$2 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=395000000000P PS=1270000U PD=1790000U
M$3 VPWR B1 \$12 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=395000000000P AD=135000000000P PS=1790000U PD=1270000U
M$4 \$12 B2 Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$5 Y B2 \$12 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$6 \$12 B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=175000000000P PS=1270000U PD=1350000U
M$7 VPWR A1 \$13 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=175000000000P AD=135000000000P PS=1350000U PD=1270000U
M$8 \$13 A2 Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$9 Y A2 \$13 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$10 \$13 A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=285000000000P PS=1270000U PD=2570000U
M$11 \$6 B1 \$3 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=169000000000P AD=87750000000P PS=1820000U PD=920000U
M$12 \$3 B2 \$6 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$13 \$6 B2 \$3 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$14 \$3 B1 \$6 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=113750000000P PS=920000U PD=1000000U
M$15 \$6 A1 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=113750000000P AD=87750000000P PS=1000000U PD=920000U
M$16 VGND A2 \$6 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=87750000000P PS=920000U PD=920000U
M$17 \$6 A2 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=87750000000P PS=920000U PD=920000U
M$18 VGND A1 \$6 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=169000000000P PS=920000U PD=1820000U
M$19 \$3 C1 Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=169000000000P
+ AD=87750000000P PS=1820000U PD=920000U
M$20 Y C1 \$3 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=169000000000P PS=920000U PD=1820000U
.ENDS sky130_fd_sc_hd__o221ai_2

.SUBCKT sky130_fd_sc_hd__a22o_2 VPB B2 B1 A1 A2 VGND X VPWR VNB
M$1 VPWR A1 \$7 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=165000000000P PS=2520000U PD=1330000U
M$2 \$7 A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=165000000000P AD=157500000000P PS=1330000U PD=1315000U
M$3 VPWR \$8 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=157500000000P AD=135000000000P PS=1315000U PD=1270000U
M$4 X \$8 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=270000000000P PS=1270000U PD=2540000U
M$5 \$8 B2 \$7 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=135000000000P PS=2520000U PD=1270000U
M$6 \$7 B1 \$8 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$7 VGND B2 \$12 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=169000000000P AD=74750000000P PS=1820000U PD=880000U
M$8 \$12 B1 \$8 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=74750000000P
+ AD=169000000000P PS=880000U PD=1820000U
M$9 \$8 A1 \$13 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=169000000000P AD=107250000000P PS=1820000U PD=980000U
M$10 \$13 A2 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=107250000000P AD=102375000000P PS=980000U PD=965000U
M$11 VGND \$8 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=102375000000P AD=87750000000P PS=965000U PD=920000U
M$12 X \$8 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=175500000000P PS=920000U PD=1840000U
.ENDS sky130_fd_sc_hd__a22o_2

.SUBCKT sky130_fd_sc_hd__dfrtp_2 VGND RESET_B Q CLK D VPWR VPB VNB
M$1 VPWR D \$5 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=109200000000P AD=65100000000P PS=1360000U PD=730000U
M$2 \$5 \$4 \$6 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=65100000000P AD=72450000000P PS=730000U PD=765000U
M$3 \$6 \$3 \$19 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=72450000000P AD=115500000000P PS=765000U PD=970000U
M$4 \$19 \$17 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=115500000000P AD=70350000000P PS=970000U PD=755000U
M$5 VPWR RESET_B \$19 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=70350000000P AD=109200000000P PS=755000U PD=1360000U
M$6 VPWR \$9 Q VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=301200000000P AD=135000000000P PS=2660000U PD=1270000U
M$7 Q \$9 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$8 \$3 CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=640000U
+ AS=166400000000P AD=86400000000P PS=1800000U PD=910000U
M$9 VPWR \$3 \$4 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=640000U
+ AS=86400000000P AD=166400000000P PS=910000U PD=1800000U
M$10 VPWR \$6 \$17 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=840000U
+ AS=218400000000P AD=129150000000P PS=2200000U PD=1185000U
M$11 \$17 \$3 \$8 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=129150000000P AD=58800000000P PS=1185000U PD=700000U
M$12 \$8 \$4 \$21 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=58800000000P AD=56700000000P PS=700000U PD=690000U
M$13 \$21 \$9 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=56700000000P AD=81900000000P PS=690000U PD=810000U
M$14 VPWR RESET_B \$9 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=81900000000P AD=56700000000P PS=810000U PD=690000U
M$15 \$9 \$8 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=56700000000P AD=113400000000P PS=690000U PD=1380000U
M$16 VGND \$9 Q VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=208700000000P AD=87750000000P PS=2020000U PD=920000U
M$17 Q \$9 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=169000000000P PS=920000U PD=1820000U
M$18 \$3 CLK VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=109200000000P AD=56700000000P PS=1360000U PD=690000U
M$19 VGND \$3 \$4 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=56700000000P AD=109200000000P PS=690000U PD=1360000U
M$20 \$6 \$3 \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=360000U
+ AS=59400000000P AD=66000000000P PS=690000U PD=745000U
M$21 \$6 \$4 \$12 VNB sky130_fd_pr__nfet_01v8 L=150000U W=360000U
+ AS=59400000000P AD=140100000000P PS=690000U PD=1100000U
M$22 \$8 \$4 \$17 VNB sky130_fd_pr__nfet_01v8 L=150000U W=360000U
+ AS=71100000000P AD=99900000000P PS=755000U PD=985000U
M$23 \$8 \$3 \$13 VNB sky130_fd_pr__nfet_01v8 L=150000U W=360000U
+ AS=71100000000P AD=66900000000P PS=755000U PD=750000U
M$24 VGND D \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=220500000000P AD=66000000000P PS=1890000U PD=745000U
M$25 \$12 \$17 \$14 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=140100000000P AD=44100000000P PS=1100000U PD=630000U
M$26 \$14 RESET_B VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=44100000000P AD=134600000000P PS=630000U PD=1150000U
M$27 \$13 \$9 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=66900000000P AD=124950000000P PS=750000U PD=1015000U
M$28 VGND RESET_B \$11 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=124950000000P AD=64050000000P PS=1015000U PD=725000U
M$29 \$11 \$8 \$9 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=64050000000P AD=109200000000P PS=725000U PD=1360000U
M$30 VGND \$6 \$17 VNB sky130_fd_pr__nfet_01v8 L=150000U W=640000U
+ AS=134600000000P AD=99900000000P PS=1150000U PD=985000U
.ENDS sky130_fd_sc_hd__dfrtp_2
