* Extracted by KLayout on : 28/07/2021 13:38

.SUBCKT DFFRAM
X$1 \$16 \$3712 \$3687 \$3743 \$1 \$16 \$153 VNB sky130_fd_sc_hd__mux2_1
X$2 \$16 \$3712 \$3306 \$3541 \$2 \$16 \$153 VNB sky130_fd_sc_hd__mux2_1
X$3 \$16 \$3270 \$3646 \$3308 \$3 \$16 \$153 VNB sky130_fd_sc_hd__mux2_1
X$4 \$16 \$3270 \$3842 \$3416 \$4 \$16 \$153 VNB sky130_fd_sc_hd__mux2_1
X$5 \$16 \$3270 \$4070 \$3311 \$5 \$16 \$153 VNB sky130_fd_sc_hd__mux2_1
X$6 \$16 \$3272 \$2794 \$3159 \$6 \$16 \$153 VNB sky130_fd_sc_hd__mux2_1
X$7 \$16 \$3272 \$4675 \$3201 \$7 \$16 \$153 VNB sky130_fd_sc_hd__mux2_1
X$8 \$153 \$8 \$398 \$9 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9 \$153 \$8 \$86 \$149 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10 \$153 \$15 \$57 \$9 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11 \$16 \$151 \$16 \$153 \$9 VNB sky130_fd_sc_hd__inv_1
X$12 \$153 \$150 \$23 \$9 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13 \$153 \$1180 \$703 \$9 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14 \$153 \$341 \$393 \$9 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15 \$153 \$312 \$549 \$9 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16 \$153 \$496 \$371 \$9 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17 \$153 \$228 \$223 \$9 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18 \$16 \$9 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19 \$16 \$9 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20 \$16 \$9 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21 \$16 \$9 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22 \$16 \$9 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23 \$16 \$9 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24 \$16 \$9 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25 \$16 \$9 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26 \$16 \$3086 \$3087 \$3088 \$10 \$16 \$153 VNB sky130_fd_sc_hd__mux2_1
X$27 \$153 \$108 \$11 \$329 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28 \$153 \$1738 \$1482 \$11 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29 \$16 \$11 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30 \$153 \$236 \$11 \$175 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31 \$153 \$719 \$11 \$600 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32 \$153 \$825 \$11 \$760 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33 \$153 \$136 \$11 \$325 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34 \$153 \$986 \$11 \$909 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35 \$153 \$107 \$11 \$20 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36 \$153 \$1025 \$11 \$1051 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37 \$153 \$1316 \$11 \$1335 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38 \$153 \$768 \$11 \$767 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39 \$153 \$36 \$11 \$176 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40 \$153 \$735 \$11 \$655 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41 \$153 \$211 \$11 \$186 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42 \$153 \$34 \$11 \$105 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43 \$153 \$875 \$11 \$1040 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44 \$153 \$718 \$11 \$641 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45 \$153 \$544 \$11 \$769 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46 \$153 \$911 \$11 \$1411 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47 \$153 \$891 \$11 \$910 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48 \$153 \$476 \$11 \$436 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49 \$153 \$1218 \$11 \$1111 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$50 \$153 \$1441 \$11 \$1410 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$51 \$153 \$1394 \$11 \$1393 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$52 \$153 \$1293 \$11 \$1199 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$53 \$153 \$153 \$11 \$1487 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$54 \$153 \$164 \$11 \$188 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$55 \$153 \$1290 \$11 \$1333 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$56 \$153 \$1288 \$11 \$1409 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$57 \$153 \$288 \$11 \$271 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$58 \$153 \$1097 \$11 \$1196 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$59 \$153 \$1506 \$11 \$1633 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$60 \$153 \$846 \$11 \$810 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$61 \$153 \$160 \$11 \$174 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$62 \$16 \$12 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$63 \$153 \$142 \$61 \$12 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$64 \$153 \$1407 \$12 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$65 \$153 \$1397 \$1254 \$12 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$66 \$153 \$198 \$267 \$12 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$67 \$153 \$219 \$189 \$12 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$68 \$153 \$579 \$425 \$12 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$69 \$153 \$722 \$670 \$12 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$70 \$153 \$408 \$407 \$12 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$71 \$153 \$1510 \$1183 \$12 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$72 \$153 \$40 \$76 \$12 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$73 \$153 \$143 \$77 \$12 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$74 \$153 \$1269 \$1268 \$12 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$75 \$153 \$437 \$422 \$12 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$76 \$153 \$45 \$62 \$12 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$77 \$153 \$118 \$81 \$12 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$78 \$153 \$1368 \$1338 \$12 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$79 \$153 \$1377 \$1185 \$12 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$80 \$153 \$1299 \$1253 \$12 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$81 \$153 \$167 \$78 \$12 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$82 \$153 \$1134 \$854 \$12 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$83 \$153 \$827 \$958 \$12 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$84 \$153 \$993 \$1026 \$12 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$85 \$153 \$992 \$826 \$12 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$86 \$153 \$1413 \$1424 \$12 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$87 \$153 \$999 \$1270 \$12 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$88 \$153 \$773 \$830 \$12 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$89 \$153 \$962 \$1043 \$12 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$90 \$153 \$828 \$1056 \$12 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$91 \$153 \$698 \$592 \$12 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$92 \$153 \$916 \$893 \$12 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$93 \$153 \$1274 \$1320 \$12 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$94 \$153 \$488 \$593 \$12 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$95 \$153 \$796 \$590 \$12 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$96 \$16 \$12 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$97 \$16 \$12 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$98 \$16 \$12 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$99 \$16 \$12 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$100 \$16 \$12 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$101 \$16 \$12 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$102 \$16 \$12 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$103 \$16 \$12 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$104 \$16 \$12 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$105 \$16 \$12 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$106 \$16 \$12 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$107 \$16 \$12 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$108 \$16 \$12 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$109 \$16 \$12 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$110 \$16 \$12 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$111 \$16 \$12 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$112 \$16 \$12 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$113 \$16 \$12 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$114 \$16 \$12 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$115 \$16 \$12 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$116 \$16 \$12 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$117 \$16 \$12 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$118 \$16 \$12 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$119 \$16 \$12 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$120 \$16 \$12 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$121 \$16 \$12 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$122 \$16 \$12 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$123 \$16 \$12 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$124 \$16 \$12 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$125 \$16 \$12 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$126 \$16 \$12 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$127 \$153 \$1406 \$13 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$128 \$153 \$699 \$593 \$13 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$129 \$153 \$220 \$81 \$13 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$130 \$153 \$882 \$893 \$13 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$131 \$153 \$147 \$62 \$13 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$132 \$153 \$41 \$78 \$13 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$133 \$153 \$1318 \$1183 \$13 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$134 \$153 \$997 \$1056 \$13 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$135 \$153 \$1114 \$1270 \$13 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$136 \$153 \$739 \$590 \$13 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$137 \$153 \$1319 \$1338 \$13 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$138 \$153 \$1226 \$1043 \$13 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$139 \$153 \$1376 \$1185 \$13 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$140 \$153 \$880 \$958 \$13 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$141 \$153 \$741 \$670 \$13 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$142 \$153 \$576 \$592 \$13 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$143 \$153 \$935 \$826 \$13 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$144 \$153 \$42 \$189 \$13 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$145 \$153 \$1369 \$1253 \$13 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$146 \$153 \$1371 \$1254 \$13 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$147 \$153 \$144 \$267 \$13 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$148 \$153 \$694 \$422 \$13 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$149 \$153 \$1133 \$854 \$13 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$150 \$153 \$934 \$1026 \$13 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$151 \$153 \$1238 \$1268 \$13 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$152 \$153 \$610 \$830 \$13 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$153 \$153 \$489 \$425 \$13 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$154 \$153 \$218 \$76 \$13 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$155 \$153 \$547 \$407 \$13 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$156 \$153 \$1448 \$1424 \$13 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$157 \$153 \$1374 \$1320 \$13 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$158 \$153 \$165 \$61 \$13 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$159 \$153 \$114 \$77 \$13 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$160 \$16 \$13 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$161 \$16 \$13 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$162 \$16 \$13 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$163 \$16 \$13 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$164 \$16 \$13 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$165 \$16 \$13 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$166 \$16 \$13 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$167 \$16 \$13 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$168 \$16 \$13 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$169 \$16 \$13 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$170 \$16 \$13 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$171 \$16 \$13 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$172 \$16 \$13 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$173 \$16 \$13 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$174 \$16 \$13 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$175 \$16 \$13 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$176 \$16 \$13 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$177 \$16 \$13 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$178 \$16 \$13 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$179 \$16 \$13 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$180 \$16 \$13 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$181 \$16 \$13 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$182 \$16 \$13 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$183 \$16 \$13 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$184 \$16 \$13 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$185 \$16 \$13 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$186 \$16 \$13 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$187 \$16 \$13 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$188 \$16 \$13 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$189 \$16 \$13 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$190 \$16 \$13 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$191 \$16 \$13 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$192 \$153 \$1539 \$14 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$193 \$153 \$1381 \$1342 \$14 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$194 \$153 \$150 \$86 \$14 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$195 \$153 \$152 \$87 \$14 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$196 \$153 \$1624 \$1568 \$14 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$197 \$153 \$1602 \$1492 \$14 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$198 \$153 \$638 \$597 \$14 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$199 \$153 \$747 \$596 \$14 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$200 \$153 \$1379 \$1278 \$14 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$201 \$153 \$805 \$762 \$14 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$202 \$153 \$806 \$706 \$14 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$203 \$153 \$148 \$85 \$14 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$204 \$153 \$746 \$761 \$14 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$205 \$153 \$1033 \$1058 \$14 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$206 \$153 \$46 \$83 \$14 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$207 \$153 \$413 \$391 \$14 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$208 \$153 \$491 \$427 \$14 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$209 \$153 \$125 \$227 \$14 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$210 \$153 \$1587 \$1340 \$14 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$211 \$153 \$226 \$84 \$14 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$212 \$153 \$647 \$676 \$14 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$213 \$153 \$170 \$50 \$14 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$214 \$153 \$171 \$277 \$14 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$215 \$153 \$809 \$836 \$14 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$216 \$153 \$1011 \$966 \$14 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$217 \$153 \$1008 \$1006 \$14 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$218 \$153 \$1009 \$943 \$14 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$219 \$153 \$1403 \$1416 \$14 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$220 \$153 \$1383 \$1302 \$14 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$221 \$153 \$1306 \$1186 \$14 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$222 \$153 \$1589 \$1565 \$14 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$223 \$153 \$1534 \$1622 \$14 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$224 \$153 \$1061 \$1147 \$14 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$225 \$16 \$14 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$226 \$16 \$14 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$227 \$16 \$14 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$228 \$16 \$14 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$229 \$16 \$14 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$230 \$16 \$14 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$231 \$16 \$14 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$232 \$16 \$14 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$233 \$16 \$14 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$234 \$16 \$14 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$235 \$16 \$14 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$236 \$16 \$14 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$237 \$16 \$14 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$238 \$16 \$14 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$239 \$16 \$14 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$240 \$16 \$14 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$241 \$16 \$14 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$242 \$16 \$14 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$243 \$16 \$14 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$244 \$16 \$14 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$245 \$16 \$14 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$246 \$16 \$14 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$247 \$16 \$14 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$248 \$16 \$14 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$249 \$16 \$14 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$250 \$16 \$14 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$251 \$16 \$14 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$252 \$16 \$14 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$253 \$16 \$14 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$254 \$16 \$14 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$255 \$16 \$14 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$256 \$16 \$14 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$257 \$153 \$15 \$86 \$63 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$258 \$153 \$10135 \$8715 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$259 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$260 \$16 \$10135 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$261 \$153 \$9878 \$9875 \$8828 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$262 \$153 \$9799 \$9875 \$9026 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$265 \$16 \$8715 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$266 \$153 \$10116 \$9831 \$8715 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$267 \$153 \$10663 \$10161 \$10006 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$268 \$153 \$10116 \$8638 \$9729 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$269 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$270 \$153 \$9604 \$9832 \$8828 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$272 \$16 \$8715 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$273 \$153 \$10012 \$9832 \$8715 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$274 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$275 \$153 \$10117 \$9879 \$9026 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$276 \$16 \$9026 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$277 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$278 \$16 \$8715 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$279 \$153 \$10136 \$10088 \$10211 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$283 \$153 \$10142 \$8638 \$9865 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$285 \$16 \$8715 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$286 \$153 \$10160 \$9765 \$8715 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$287 \$153 \$10090 \$9765 \$8828 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$288 \$16 \$8828 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$289 \$153 \$10091 \$8638 \$9866 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$291 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$292 \$16 \$9026 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$293 \$153 \$10118 \$9793 \$8828 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$294 \$16 \$8828 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$296 \$16 \$6666 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$297 \$153 \$6666 \$10143 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$299 \$153 \$9966 \$8726 \$9836 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$301 \$153 \$9946 \$9880 \$8436 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$302 \$16 \$10226 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$304 \$153 \$8839 \$8436 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$306 \$153 \$10017 \$9838 \$8436 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$308 \$153 \$9227 \$9026 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$309 \$153 \$10119 \$8340 \$8638 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$310 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$311 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$312 \$153 \$10120 \$8340 \$10088 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$314 \$153 \$10036 \$3910 \$10093 \$10144 \$10145 \$9075 \$10007 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$315 \$153 \$10036 \$3687 \$9967 \$10146 \$10147 \$8955 \$10007 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$316 \$16 \$7934 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$318 \$153 \$10095 \$8614 \$9868 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$319 \$16 \$8647 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$321 \$153 \$10162 \$9900 \$8816 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$322 \$153 \$10148 \$8789 \$9868 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$323 \$16 \$8816 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$324 \$153 \$10121 \$9794 \$8816 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$325 \$153 \$10121 \$8804 \$9902 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$326 \$16 \$8816 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$329 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$331 \$153 \$10163 \$9795 \$8816 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$332 \$153 \$10149 \$8789 \$9720 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$333 \$153 \$10064 \$8727 \$9720 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$334 \$153 \$10137 \$8277 \$9720 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$335 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$337 \$153 \$10150 \$8804 \$9842 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$338 \$153 \$10164 \$9811 \$8816 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$339 \$153 \$10038 \$8277 \$9842 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$340 \$153 \$10066 \$8651 \$9586 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$341 \$16 \$8816 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$342 \$16 \$8441 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$343 \$153 \$10039 \$8727 \$9815 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$346 \$16 \$5765 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$347 \$16 \$10165 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$348 \$16 \$10166 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$350 \$153 \$10096 \$9884 \$8890 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$351 \$16 \$7949 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$352 \$16 \$7949 \$16 \$153 \$10167 VNB sky130_fd_sc_hd__clkbuf_2
X$353 \$153 \$10167 \$4668 \$8697 \$10151 \$10122 \$10152 \$10082 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$354 \$16 \$8890 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$355 \$16 \$8697 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$358 \$16 \$10122 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$359 \$16 \$10180 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$360 \$153 \$10205 \$8886 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$361 \$153 \$10139 \$8816 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$362 \$16 \$10139 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$363 \$153 \$9690 \$8610 \$9746 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$366 \$153 \$10238 \$8728 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$368 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$369 \$153 \$10123 \$8340 \$10098 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$370 \$153 \$10138 \$8340 \$9133 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$373 \$153 \$9817 \$8818 \$9845 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$375 \$153 \$9970 \$8340 \$9174 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$376 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$377 \$16 \$10247 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$378 \$16 \$8789 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$379 \$16 \$8277 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$380 \$153 \$10168 \$10021 \$9214 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$381 \$16 \$9214 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$382 \$16 \$9047 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$383 \$16 \$9031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$385 \$153 \$10124 \$10021 \$9031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$386 \$16 \$9174 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$388 \$16 \$9045 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$389 \$153 \$9951 \$10000 \$9045 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$390 \$153 \$10124 \$9133 \$10216 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$392 \$153 \$10102 \$8842 \$9871 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$394 \$16 \$8820 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$395 \$16 \$8313 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$397 \$16 \$9045 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$398 \$153 \$10169 \$10083 \$9045 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$400 \$16 \$7996 \$16 \$153 \$9953 VNB sky130_fd_sc_hd__inv_1
X$401 \$16 \$8936 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$403 \$153 \$10170 \$10083 \$9031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$404 \$153 \$10070 \$8842 \$9953 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$407 \$153 \$10103 \$9934 \$9045 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$408 \$153 \$10171 \$9934 \$9188 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$409 \$153 \$10172 \$10022 \$9045 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$410 \$16 \$9253 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$411 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$412 \$16 \$8624 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$415 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$417 \$153 \$10155 \$9252 \$10009 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$418 \$153 \$10156 \$9047 \$10009 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$420 \$153 \$10072 \$8676 \$10104 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$421 \$153 \$10125 \$10024 \$9031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$422 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$425 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$426 \$16 \$9045 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$427 \$153 \$9890 \$10157 \$9045 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$429 \$153 \$10105 \$8842 \$9872 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$430 \$153 \$9937 \$10157 \$9031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$431 \$16 \$9045 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$432 \$16 \$7949 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$433 \$16 \$7949 \$16 \$153 \$10075 VNB sky130_fd_sc_hd__clkbuf_2
X$435 \$153 \$10126 \$10010 \$9045 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$437 \$16 \$10101 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$438 \$153 \$10173 \$10010 \$9031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$439 \$153 \$10075 \$4262 \$10045 \$10101 \$10158 \$10127 \$10220 \$16 \$16
+ VNB sky130_fd_sc_hd__mux4_1
X$441 \$153 \$10075 \$4141 \$10044 \$10123 \$10159 \$9856 \$10220 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$442 \$153 \$10174 \$8340 \$9103 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$443 \$153 \$10127 \$8340 \$9256 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$444 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$447 \$153 \$10128 \$9913 \$9154 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$448 \$153 \$10128 \$9103 \$9981 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$449 \$153 \$10140 \$9940 \$9154 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$450 \$153 \$10140 \$9103 \$10108 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$451 \$16 \$8879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$453 \$16 \$9134 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$455 \$153 \$10129 \$9940 \$9134 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$457 \$16 \$9154 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$458 \$153 \$10130 \$10025 \$9154 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$459 \$153 \$9958 \$10025 \$8927 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$460 \$16 \$8927 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$461 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$464 \$16 \$8927 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$465 \$153 \$10175 \$10085 \$8927 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$466 \$153 \$10175 \$9256 \$10110 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$467 \$153 \$10131 \$10085 \$9035 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$468 \$153 \$10131 \$8977 \$10110 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$469 \$16 \$8879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$471 \$153 \$10027 \$10111 \$8893 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$472 \$16 \$8893 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$474 \$153 \$10132 \$10111 \$8927 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$475 \$153 \$10132 \$9256 \$9988 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$477 \$16 \$7076 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$478 \$153 \$10133 \$9256 \$10112 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$480 \$16 \$8453 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$481 \$16 \$9034 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$482 \$153 \$10141 \$8923 \$9961 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$483 \$153 \$10182 \$9059 \$9961 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$485 \$153 \$10133 \$10028 \$8927 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$486 \$153 \$10113 \$9103 \$10112 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$487 \$16 \$8893 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$488 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$490 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$491 \$16 \$8927 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$492 \$153 \$10177 \$9991 \$8927 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$494 \$153 \$10134 \$9103 \$10005 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$495 \$153 \$10134 \$9991 \$9154 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$496 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$499 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$500 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$501 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$502 \$153 \$6708 \$10135 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$503 \$16 \$6708 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$504 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$506 \$153 \$10206 \$10303 \$10006 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$508 \$16 \$8828 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$509 \$153 \$10207 \$10330 \$10006 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$510 \$153 \$10208 \$10088 \$10245 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$511 \$153 \$9945 \$9831 \$9026 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$512 \$153 \$10183 \$10705 \$10006 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$514 \$16 \$9026 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$515 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$516 \$153 \$10209 \$10303 \$10210 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$518 \$153 \$10184 \$9832 \$9026 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$519 \$16 \$8828 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$520 \$16 \$9026 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$522 \$153 \$10296 \$10276 \$10211 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$523 \$153 \$10227 \$10161 \$10211 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$525 \$153 \$10178 \$9879 \$8436 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$527 \$153 \$10142 \$9879 \$8715 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$528 \$16 \$8436 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$529 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$531 \$153 \$10185 \$9765 \$9026 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$533 \$153 \$10160 \$8638 \$9740 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$534 \$153 \$10185 \$8726 \$9740 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$536 \$153 \$10186 \$10199 \$10200 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$538 \$153 \$10213 \$10303 \$10212 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$539 \$153 \$10187 \$10161 \$10212 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$540 \$16 \$10200 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$542 \$153 \$10118 \$8885 \$9866 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$544 \$153 \$10143 \$8828 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$545 \$16 \$10295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$546 \$16 \$10200 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$547 \$16 \$6646 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$548 \$153 \$6646 \$8839 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$550 \$16 \$8436 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$551 \$16 \$6820 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$552 \$153 \$6820 \$9227 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$553 \$153 \$6722 \$10042 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$554 \$153 \$9741 \$8209 \$9567 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$556 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$558 \$153 \$10230 \$8340 \$8726 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$559 \$16 \$10088 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$560 \$153 \$10036 \$3911 \$10094 \$10201 \$10202 \$8787 \$10007 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$561 \$16 \$9336 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$562 \$16 \$8787 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$563 \$16 \$8957 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$564 \$16 \$9075 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$565 \$153 \$10188 \$8727 \$9868 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$567 \$16 \$7934 \$16 \$153 \$10007 VNB sky130_fd_sc_hd__clkbuf_2
X$569 \$153 \$10188 \$9900 \$8886 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$570 \$16 \$8886 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$572 \$153 \$10148 \$9900 \$8898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$573 \$16 \$8898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$574 \$16 \$8806 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$575 \$16 \$10080 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$577 \$153 \$10214 \$8277 \$9902 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$579 \$153 \$10189 \$9794 \$8898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$580 \$153 \$10189 \$8789 \$9902 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$581 \$16 \$8898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$582 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$583 \$153 \$10149 \$9795 \$8898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$584 \$16 \$8898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$585 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$588 \$16 \$6669 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$589 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$590 \$153 \$10190 \$9796 \$8898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$591 \$153 \$10190 \$8789 \$9842 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$592 \$16 \$8898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$593 \$16 \$8898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$594 \$153 \$10191 \$9811 \$8898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$596 \$16 \$10215 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$597 \$16 \$10179 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$599 \$153 \$10191 \$8789 \$9586 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$600 \$153 \$10167 \$3978 \$8441 \$10179 \$9885 \$10203 \$10082 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$602 \$16 \$5765 \$16 \$153 \$9550 VNB sky130_fd_sc_hd__clkbuf_2
X$603 \$153 \$10167 \$3400 \$8634 \$10166 \$10180 \$10040 \$10082 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$605 \$153 \$10167 \$4070 \$8487 \$10357 \$10181 \$10138 \$10082 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$606 \$153 \$10310 \$8277 \$9586 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$607 \$16 \$10181 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$608 \$16 \$9845 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$609 \$16 \$8727 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$610 \$153 \$10097 \$8686 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$612 \$153 \$10067 \$8789 \$9845 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$614 \$153 \$10408 \$8898 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$615 \$153 \$10192 \$8340 \$8804 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$616 \$153 \$9906 \$8789 \$9746 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$619 \$153 \$10154 \$8340 \$10401 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$620 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$621 \$153 \$10203 \$8340 \$8842 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$622 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$623 \$153 \$10152 \$8340 \$8917 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$624 \$16 \$8839 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$625 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$627 \$153 \$10081 \$8340 \$9252 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$628 \$153 \$9972 \$9278 \$9453 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$629 \$153 \$10168 \$9047 \$10216 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$630 \$16 \$9188 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$631 \$16 \$8842 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$632 \$16 \$9188 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$633 \$153 \$10231 \$10000 \$9188 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$635 \$153 \$10099 \$9174 \$10216 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$636 \$16 \$8719 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$637 \$16 \$9031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$638 \$153 \$10193 \$10000 \$9031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$639 \$153 \$10217 \$9278 \$9871 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$640 \$153 \$10193 \$9133 \$9871 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$641 \$153 \$10169 \$9174 \$9953 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$643 \$153 \$10218 \$9047 \$9953 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$644 \$16 \$9031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$645 \$16 \$7996 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$646 \$153 \$10170 \$9133 \$9953 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$647 \$16 \$9045 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$648 \$16 \$9214 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$649 \$153 \$10194 \$9934 \$9214 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$650 \$153 \$10194 \$9047 \$9927 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$651 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$654 \$153 \$10171 \$8917 \$9927 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$655 \$16 \$9045 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$656 \$153 \$10172 \$9174 \$10009 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$657 \$153 \$10155 \$10022 \$9253 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$658 \$16 \$9253 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$659 \$16 \$9188 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$660 \$153 \$10235 \$10024 \$9188 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$663 \$16 \$9214 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$665 \$16 \$9275 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$666 \$153 \$10195 \$10024 \$9275 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$667 \$153 \$10195 \$9278 \$10104 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$669 \$16 \$8807 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$670 \$153 \$9891 \$10157 \$8807 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$671 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$673 \$153 \$10219 \$9252 \$9872 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$674 \$16 \$8704 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$675 \$16 \$9188 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$676 \$153 \$10196 \$9047 \$9872 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$677 \$153 \$10106 \$10010 \$9188 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$678 \$153 \$10236 \$9252 \$9955 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$679 \$153 \$10237 \$9047 \$9955 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$681 \$16 \$7934 \$16 \$153 \$10220 VNB sky130_fd_sc_hd__clkbuf_2
X$682 \$16 \$7934 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$684 \$153 \$10221 \$9278 \$9955 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$685 \$153 \$10173 \$9133 \$9955 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$686 \$16 \$10154 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$687 \$153 \$10075 \$2960 \$10069 \$10154 \$10204 \$10049 \$10220 \$16 \$16
+ VNB sky130_fd_sc_hd__mux4_1
X$688 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$689 \$16 \$10069 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$690 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$692 \$16 \$8313 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$693 \$16 \$9103 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$694 \$16 \$10238 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$695 \$153 \$10107 \$9256 \$9981 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$696 \$153 \$10238 \$8927 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$698 \$153 \$10139 \$9154 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$700 \$153 \$10239 \$9940 \$8879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$701 \$16 \$10139 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$702 \$16 \$10205 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$704 \$16 \$9035 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$705 \$153 \$10197 \$9940 \$9035 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$706 \$153 \$10197 \$8977 \$10108 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$707 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$708 \$16 \$9035 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$710 \$153 \$10109 \$10025 \$9035 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$711 \$153 \$10240 \$10025 \$8879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$712 \$16 \$10097 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$713 \$16 \$8879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$714 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$715 \$153 \$10198 \$10085 \$8879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$717 \$153 \$10198 \$8923 \$10110 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$718 \$16 \$8879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$719 \$16 \$8702 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$720 \$16 \$8624 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$721 \$153 \$10176 \$9256 \$10222 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$722 \$153 \$10242 \$10111 \$8879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$723 \$153 \$10243 \$10111 \$9134 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$725 \$16 \$9134 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$727 \$153 \$10223 \$8977 \$9988 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$729 \$16 \$8879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$730 \$153 \$10141 \$9860 \$8879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$731 \$153 \$10182 \$9860 \$9034 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$732 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$734 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$736 \$153 \$10224 \$8977 \$10112 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$737 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$739 \$153 \$10054 \$8965 \$10112 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$740 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$741 \$16 \$8879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$743 \$153 \$10177 \$9256 \$10005 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$744 \$153 \$10115 \$8996 \$10005 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$746 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$747 \$16 \$9035 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$748 \$153 \$10244 \$9991 \$9035 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$749 \$153 \$8714 \$7462 \$8777 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$750 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$751 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$752 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$753 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$755 \$153 \$11884 \$11733 \$10368 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$756 \$16 \$10368 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$758 \$153 \$11854 \$11733 \$10367 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$759 \$153 \$11854 \$10330 \$11717 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$761 \$16 \$11757 \$11347 \$11885 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$762 \$153 \$11870 \$10161 \$11717 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$764 \$153 \$11886 \$11751 \$10368 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$765 \$16 \$10368 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$766 \$16 \$11757 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$767 \$16 \$10348 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$768 \$16 \$11898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$769 \$153 \$11812 \$11751 \$10367 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$772 \$16 \$11898 \$16 \$153 \$11718 VNB sky130_fd_sc_hd__inv_1
X$773 \$153 \$11887 \$11631 \$10226 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$774 \$153 \$11855 \$11631 \$10367 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$775 \$153 \$11855 \$10330 \$11650 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$776 \$153 \$11871 \$10088 \$11650 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$777 \$16 \$11888 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$780 \$16 \$12013 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$781 \$16 \$11721 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$782 \$153 \$11889 \$11632 \$10368 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$783 \$153 \$11890 \$11632 \$10367 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$784 \$16 \$11721 \$16 \$153 \$11560 VNB sky130_fd_sc_hd__inv_1
X$785 \$153 \$11891 \$11633 \$10368 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$788 \$153 \$11890 \$10330 \$11560 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$789 \$153 \$11892 \$11633 \$10226 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$790 \$16 \$11800 \$16 \$153 \$11652 VNB sky130_fd_sc_hd__inv_1
X$791 \$16 \$10226 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$792 \$16 \$10367 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$793 \$153 \$11893 \$11735 \$10367 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$794 \$16 \$10476 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$795 \$16 \$11800 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$796 \$16 \$11800 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$799 \$153 \$11813 \$11735 \$10368 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$800 \$16 \$11795 \$16 \$153 \$11719 VNB sky130_fd_sc_hd__inv_1
X$802 \$153 \$11894 \$11801 \$10367 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$803 \$153 \$11894 \$10330 \$11655 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$804 \$153 \$11834 \$10705 \$11655 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$805 \$16 \$10200 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$807 \$153 \$11896 \$11801 \$10368 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$808 \$153 \$11895 \$10161 \$11655 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$810 \$16 \$11805 \$11856 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$811 \$16 \$11690 \$16 \$153 \$11594 VNB sky130_fd_sc_hd__clkbuf_2
X$812 \$16 \$11760 \$16 \$153 \$11814 VNB sky130_fd_sc_hd__clkbuf_2
X$813 \$16 \$11944 \$10888 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$814 \$16 \$11944 \$10890 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$815 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$816 \$16 \$11736 \$16 \$153 \$11636 VNB sky130_fd_sc_hd__clkbuf_2
X$817 \$16 \$11805 \$11897 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$818 \$16 \$11836 \$16 \$153 \$11898 VNB sky130_fd_sc_hd__clkbuf_2
X$820 \$16 \$11816 \$16 \$153 \$11794 VNB sky130_fd_sc_hd__clkbuf_2
X$822 \$16 \$11898 \$11275 \$11899 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$823 \$16 \$11835 \$16 \$153 \$11757 VNB sky130_fd_sc_hd__clkbuf_2
X$824 \$16 \$11898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$825 \$153 \$11817 \$11737 \$10514 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$826 \$153 \$11819 \$11737 \$10605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$827 \$16 \$10605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$829 \$16 \$11987 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$830 \$16 \$10526 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$832 \$153 \$11820 \$11737 \$10382 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$833 \$153 \$11872 \$10344 \$11818 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$834 \$16 \$10382 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$835 \$153 \$11618 \$10247 \$11838 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$836 \$153 \$11873 \$10516 \$11838 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$837 \$16 \$10526 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$838 \$16 \$11794 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$839 \$16 \$11888 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$840 \$16 \$11721 \$11275 \$11900 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$843 \$16 \$10514 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$844 \$153 \$11619 \$10098 \$11838 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$845 \$16 \$10606 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$846 \$16 \$12013 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$847 \$153 \$11901 \$11658 \$10514 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$848 \$153 \$11874 \$10516 \$11562 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$849 \$153 \$11901 \$10538 \$11562 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$851 \$16 \$10382 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$852 \$16 \$11721 \$16 \$153 \$11660 VNB sky130_fd_sc_hd__inv_1
X$854 \$153 \$11875 \$10344 \$11562 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$856 \$153 \$11876 \$10516 \$11660 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$858 \$153 \$11857 \$11967 \$10514 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$859 \$153 \$11857 \$10538 \$11660 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$860 \$153 \$11877 \$10344 \$11660 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$861 \$16 \$11995 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$863 \$153 \$11738 \$11639 \$10514 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$864 \$16 \$10514 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$866 \$153 \$11902 \$11639 \$10526 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$867 \$16 \$11795 \$11164 \$11903 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$868 \$153 \$11905 \$11739 \$10526 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$870 \$16 \$11795 \$16 \$153 \$11563 VNB sky130_fd_sc_hd__inv_1
X$871 \$153 \$11878 \$12174 \$11869 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$872 \$153 \$11905 \$10516 \$11563 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$873 \$153 \$11879 \$10538 \$11563 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$875 \$16 \$10298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$876 \$16 \$10514 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$877 \$153 \$11373 \$11806 \$10382 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$879 \$16 \$11814 \$16 \$153 \$11906 VNB sky130_fd_sc_hd__inv_1
X$882 \$153 \$11904 \$10686 \$11488 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$883 \$16 \$8734 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$884 \$153 \$11907 \$11806 \$10526 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$885 \$16 \$10526 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$886 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$887 \$153 \$8540 \$8340 \$12476 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$888 \$153 \$11767 \$10686 \$11564 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$890 \$153 \$11770 \$11741 \$10809 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$891 \$16 \$10809 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$893 \$153 \$11823 \$11741 \$10551 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$894 \$153 \$11908 \$11741 \$10386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$895 \$16 \$10551 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$896 \$16 \$10551 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$899 \$153 \$11769 \$10833 \$11724 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$900 \$153 \$11909 \$11641 \$10473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$902 \$16 \$10551 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$903 \$153 \$11858 \$11666 \$10551 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$904 \$153 \$11909 \$10501 \$11665 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$905 \$16 \$10735 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$908 \$153 \$11858 \$10471 \$11513 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$910 \$16 \$10300 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$911 \$16 \$10735 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$912 \$153 \$11859 \$11742 \$10735 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$913 \$153 \$11859 \$10919 \$11669 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$915 \$153 \$11910 \$11880 \$10473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$917 \$153 \$11929 \$10714 \$11669 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$918 \$16 \$10611 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$919 \$153 \$11744 \$11880 \$10611 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$920 \$16 \$11627 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$921 \$16 \$11412 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$922 \$16 \$10300 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$923 \$153 \$11911 \$11807 \$10300 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$924 \$16 \$10809 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$925 \$16 \$11627 \$11412 \$11912 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$928 \$16 \$10578 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$929 \$153 \$11860 \$11807 \$10809 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$930 \$153 \$11860 \$10714 \$11954 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$932 \$153 \$11861 \$11645 \$10809 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$933 \$153 \$11861 \$10714 \$11727 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$934 \$16 \$11412 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$936 \$153 \$11624 \$10833 \$11727 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$937 \$16 \$11798 \$11412 \$11913 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$939 \$16 \$11483 \$11412 \$11914 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$940 \$153 \$11862 \$11808 \$10473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$941 \$153 \$11863 \$10472 \$11825 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$942 \$153 \$11862 \$10501 \$11825 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$943 \$16 \$10551 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$945 \$153 \$11864 \$11808 \$10551 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$946 \$153 \$11864 \$10471 \$11825 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$947 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$949 \$16 \$11546 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$950 \$153 \$11748 \$11780 \$11803 \$11781 \$11782 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$951 \$153 \$11780 \$11782 \$11915 \$11781 \$11803 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$952 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$954 \$16 \$11846 \$16 \$153 \$11214 VNB sky130_fd_sc_hd__clkbuf_2
X$955 \$16 \$11847 \$16 \$153 \$11496 VNB sky130_fd_sc_hd__clkbuf_2
X$957 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$958 \$16 \$11783 \$16 \$153 \$11627 VNB sky130_fd_sc_hd__clkbuf_2
X$959 \$153 \$8675 \$8340 \$11881 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$960 \$153 \$11865 \$11809 \$10564 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$961 \$153 \$11865 \$10642 \$11827 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$963 \$16 \$11824 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$965 \$16 \$11930 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$966 \$153 \$11828 \$11809 \$10446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$967 \$16 \$10346 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$968 \$16 \$10446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$969 \$16 \$12009 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$970 \$16 \$10564 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$971 \$153 \$11866 \$11628 \$10564 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$972 \$153 \$11866 \$10642 \$11829 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$976 \$16 \$11772 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$977 \$153 \$11882 \$10587 \$11829 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$978 \$16 \$11930 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$979 \$16 \$10617 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$980 \$153 \$11916 \$11629 \$10617 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$981 \$153 \$11917 \$11629 \$10446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$982 \$16 \$10446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$983 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$984 \$16 \$10467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$986 \$153 \$11918 \$11709 \$10467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$987 \$16 \$10617 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$988 \$153 \$11919 \$11709 \$10617 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$989 \$153 \$11920 \$11709 \$10392 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$990 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$991 \$16 \$11945 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$993 \$16 \$10564 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$994 \$153 \$11867 \$11681 \$10564 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$995 \$153 \$11867 \$10642 \$11730 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$997 \$153 \$11922 \$11587 \$10467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$998 \$153 \$11922 \$10587 \$11731 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$999 \$16 \$10564 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1002 \$16 \$11459 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1003 \$153 \$11883 \$10642 \$11731 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1005 \$16 \$10392 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1006 \$16 \$11798 \$11229 \$11924 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$1007 \$153 \$11923 \$11588 \$10392 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1008 \$16 \$11627 \$16 \$153 \$13451 VNB sky130_fd_sc_hd__inv_1
X$1009 \$16 \$10564 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1010 \$153 \$11925 \$11588 \$10564 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1013 \$16 \$10564 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1014 \$16 \$11798 \$16 \$153 \$11926 VNB sky130_fd_sc_hd__inv_1
X$1015 \$153 \$11927 \$11648 \$10564 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1016 \$16 \$11390 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1017 \$16 \$11798 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1018 \$16 \$10617 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1019 \$153 \$11928 \$11648 \$10617 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1020 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$1021 \$153 \$11154 \$10815 \$11022 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1023 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$1024 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$1025 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$1026 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$1027 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$1029 \$153 \$11884 \$10303 \$11717 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1031 \$153 \$11959 \$11733 \$10200 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1032 \$16 \$10200 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1033 \$16 \$10367 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1035 \$153 \$11870 \$11733 \$10226 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1036 \$16 \$11757 \$16 \$153 \$11717 VNB sky130_fd_sc_hd__inv_1
X$1037 \$153 \$11960 \$11751 \$10200 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1039 \$16 \$10200 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1040 \$153 \$11886 \$10303 \$11718 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1042 \$16 \$11949 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1043 \$153 \$11751 \$11949 \$12056 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$1044 \$16 \$10367 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1046 \$153 \$11871 \$11631 \$10200 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1047 \$153 \$11887 \$10161 \$11650 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1049 \$16 \$11794 \$11347 \$11931 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$1050 \$153 \$11631 \$11888 \$11931 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$1051 \$16 \$11721 \$11347 \$11961 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$1052 \$153 \$11932 \$11632 \$10226 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1053 \$153 \$11932 \$10161 \$11560 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1054 \$16 \$10368 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1055 \$16 \$10226 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1056 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$1058 \$153 \$11889 \$10303 \$11560 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1059 \$16 \$10367 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1060 \$153 \$11933 \$11633 \$10367 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1061 \$153 \$11891 \$10303 \$11652 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1062 \$153 \$11633 \$11897 \$11934 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$1063 \$16 \$11800 \$11238 \$11934 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$1066 \$16 \$10555 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1068 \$153 \$11962 \$11735 \$10226 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1069 \$153 \$11893 \$10330 \$11719 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1070 \$153 \$11962 \$10161 \$11719 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1071 \$153 \$11735 \$11995 \$11935 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$1072 \$16 \$11795 \$11238 \$11935 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$1074 \$153 \$11895 \$11801 \$10226 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1075 \$16 \$10226 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1076 \$153 \$11963 \$11801 \$10200 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1077 \$153 \$11896 \$10303 \$11655 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1078 \$16 \$11943 \$16 \$153 \$11994 VNB sky130_fd_sc_hd__clkbuf_2
X$1079 \$16 \$8340 \$16 \$153 \$11943 VNB sky130_fd_sc_hd__clkbuf_2
X$1080 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1081 \$16 \$11944 \$11114 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$1083 \$16 \$11943 \$16 \$153 \$11944 VNB sky130_fd_sc_hd__clkbuf_2
X$1084 \$16 \$11943 \$16 \$153 \$11805 VNB sky130_fd_sc_hd__clkbuf_2
X$1085 \$16 \$11944 \$10523 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$1086 \$16 \$11944 \$10522 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$1087 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1088 \$153 \$10321 \$8340 \$12057 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1089 \$153 \$11737 \$11949 \$11899 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$1090 \$16 \$12057 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1091 \$16 \$11949 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1092 \$16 \$10348 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1093 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$1095 \$16 \$11898 \$16 \$153 \$11818 VNB sky130_fd_sc_hd__inv_1
X$1096 \$16 \$10514 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1097 \$16 \$11898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1099 \$153 \$11964 \$11737 \$10526 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1100 \$153 \$11872 \$11737 \$10606 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1101 \$153 \$11657 \$11987 \$11965 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$1104 \$153 \$11873 \$11657 \$10526 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1105 \$153 \$11936 \$11657 \$10606 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1106 \$153 \$11658 \$11888 \$11966 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$1107 \$153 \$11936 \$10344 \$11838 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1110 \$16 \$11794 \$16 \$153 \$11562 VNB sky130_fd_sc_hd__inv_1
X$1111 \$16 \$11794 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1112 \$16 \$10744 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1113 \$153 \$11875 \$11658 \$10606 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1114 \$16 \$10606 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1115 \$153 \$11876 \$11967 \$10526 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1116 \$153 \$11950 \$10686 \$11562 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1118 \$16 \$11800 \$11164 \$11951 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$1120 \$16 \$10526 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1122 \$153 \$11639 \$11897 \$11951 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$1123 \$153 \$11904 \$11639 \$10605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1124 \$153 \$11968 \$11639 \$10606 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1125 \$16 \$10606 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1126 \$16 \$10413 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1128 \$16 \$10706 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1130 \$153 \$11739 \$11995 \$11903 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$1132 \$153 \$11821 \$11739 \$10605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1134 \$153 \$11879 \$11739 \$10514 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1135 \$16 \$10514 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1136 \$16 \$11814 \$11164 \$11969 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$1139 \$153 \$11952 \$10344 \$11563 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1140 \$153 \$11953 \$11806 \$10514 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1141 \$153 \$11970 \$11806 \$10606 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1142 \$153 \$11953 \$10538 \$11906 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1143 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1144 \$16 \$10606 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1145 \$16 \$10605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1147 \$153 \$11907 \$10516 \$11906 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1149 \$16 \$12068 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1150 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1151 \$153 \$8767 \$8340 \$12068 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1153 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1154 \$153 \$9886 \$8340 \$12217 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1155 \$16 \$10611 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1156 \$16 \$12309 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1158 \$16 \$10578 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1160 \$153 \$11971 \$11741 \$10578 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1162 \$153 \$11972 \$11641 \$10551 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1163 \$153 \$11908 \$10472 \$11724 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1164 \$153 \$11972 \$10471 \$11665 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1165 \$16 \$12165 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1167 \$16 \$10473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1169 \$153 \$11973 \$11666 \$10473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1170 \$16 \$11772 \$11378 \$11974 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$1171 \$153 \$11667 \$11666 \$10735 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1172 \$16 \$11772 \$16 \$153 \$11513 VNB sky130_fd_sc_hd__inv_1
X$1173 \$153 \$11975 \$11742 \$10386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1175 \$153 \$11929 \$11742 \$10809 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1176 \$153 \$11937 \$11880 \$10809 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1177 \$153 \$11937 \$10714 \$11725 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1178 \$153 \$11910 \$10501 \$11725 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1180 \$16 \$11945 \$16 \$153 \$11725 VNB sky130_fd_sc_hd__inv_1
X$1181 \$16 \$11945 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1183 \$16 \$11945 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1185 \$16 \$10386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1186 \$153 \$11976 \$11807 \$10386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1187 \$153 \$11844 \$10919 \$11954 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1188 \$153 \$11938 \$11807 \$10578 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1189 \$153 \$11938 \$10370 \$11954 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1191 \$153 \$11977 \$11645 \$10300 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1192 \$16 \$10300 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1193 \$16 \$10649 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1194 \$16 \$10578 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1195 \$153 \$11978 \$11645 \$10578 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1196 \$153 \$11645 \$11921 \$11913 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$1197 \$16 \$10473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1198 \$16 \$11483 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1200 \$153 \$11808 \$11946 \$11914 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$1202 \$16 \$10735 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1203 \$153 \$11939 \$11808 \$10735 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1204 \$153 \$11939 \$10919 \$11825 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1205 \$153 \$11955 \$10714 \$11825 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1206 \$16 \$11483 \$16 \$153 \$11825 VNB sky130_fd_sc_hd__inv_1
X$1207 \$16 \$11483 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1209 \$16 \$11956 \$16 \$153 \$11930 VNB sky130_fd_sc_hd__clkbuf_2
X$1210 \$153 \$11979 \$11781 \$11803 \$11780 \$11782 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$1211 \$153 \$11956 \$11782 \$11803 \$11781 \$11780 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$1212 \$16 \$11947 \$16 \$153 \$12032 VNB sky130_fd_sc_hd__clkbuf_2
X$1213 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1214 \$153 \$7833 \$8340 \$12182 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1215 \$16 \$11848 \$16 \$153 \$11798 VNB sky130_fd_sc_hd__clkbuf_2
X$1216 \$16 \$12182 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1217 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$1220 \$16 \$11881 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1222 \$153 \$11948 \$11809 \$10467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1223 \$153 \$11948 \$10587 \$11827 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1224 \$16 \$10467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1225 \$153 \$11940 \$11809 \$10617 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1226 \$16 \$10617 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1228 \$16 \$11772 \$11504 \$11980 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$1230 \$153 \$11940 \$10560 \$11827 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1231 \$16 \$10617 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1232 \$16 \$11772 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1233 \$16 \$10467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1234 \$153 \$11882 \$11628 \$10467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1235 \$16 \$11772 \$16 \$153 \$11829 VNB sky130_fd_sc_hd__inv_1
X$1237 \$16 \$10392 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1238 \$153 \$11981 \$11629 \$10392 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1239 \$16 \$11930 \$16 \$153 \$11678 VNB sky130_fd_sc_hd__inv_1
X$1241 \$16 \$12032 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1242 \$16 \$10467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1243 \$153 \$11850 \$11629 \$10467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1245 \$16 \$10564 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1246 \$153 \$11941 \$11709 \$10564 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1247 \$153 \$11941 \$10642 \$11680 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1248 \$16 \$12032 \$16 \$153 \$11680 VNB sky130_fd_sc_hd__inv_1
X$1249 \$16 \$12032 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1250 \$16 \$10736 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1254 \$16 \$10467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1255 \$153 \$11919 \$10560 \$11680 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1256 \$153 \$11982 \$11681 \$10467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1257 \$16 \$11945 \$16 \$153 \$11730 VNB sky130_fd_sc_hd__inv_1
X$1258 \$16 \$11983 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1259 \$153 \$11984 \$11681 \$10617 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1260 \$16 \$10617 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1262 \$16 \$11921 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1263 \$16 \$10392 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1265 \$153 \$11831 \$11587 \$10392 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1266 \$153 \$11883 \$11587 \$10564 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1267 \$153 \$11851 \$10560 \$11731 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1269 \$153 \$11648 \$11921 \$11924 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$1271 \$153 \$11957 \$11942 \$11958 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1273 \$153 \$11985 \$11588 \$10617 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1274 \$153 \$11460 \$10694 \$11390 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1275 \$153 \$11319 \$10285 \$11390 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1276 \$153 \$11261 \$10376 \$11390 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1278 \$16 \$10392 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1280 \$153 \$11986 \$11648 \$10392 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1281 \$153 \$10425 \$10376 \$10801 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1282 \$153 \$10452 \$10587 \$10801 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1283 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$1284 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$1285 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$1286 \$153 \$7393 \$6794 \$6855 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1287 \$153 \$7465 \$6996 \$7552 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1289 \$153 \$7499 \$7319 \$6860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1290 \$153 \$7019 \$6732 \$7078 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1291 \$16 \$6860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1293 \$16 \$6915 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1294 \$153 \$7247 \$6995 \$7078 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1295 \$16 \$6792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1296 \$153 \$7319 \$7333 \$7434 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$1297 \$153 \$7053 \$7547 \$7394 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$1298 \$16 \$7378 \$7233 \$7434 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$1300 \$153 \$7281 \$6930 \$7137 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1302 \$16 \$7381 \$16 \$153 \$7137 VNB sky130_fd_sc_hd__inv_1
X$1303 \$16 \$6783 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1305 \$153 \$7500 \$7320 \$6907 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1306 \$16 \$6907 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1307 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$1308 \$153 \$7435 \$7320 \$6783 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1309 \$153 \$7435 \$6749 \$7140 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1312 \$153 \$7501 \$7234 \$6860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1313 \$153 \$7396 \$6930 \$7141 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1314 \$153 \$7397 \$6996 \$7141 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1316 \$16 \$7466 \$16 \$153 \$7141 VNB sky130_fd_sc_hd__inv_1
X$1317 \$16 \$7467 \$16 \$153 \$7158 VNB sky130_fd_sc_hd__clkbuf_2
X$1318 \$153 \$7234 \$7335 \$7468 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$1320 \$153 \$7436 \$7235 \$6860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1321 \$153 \$7436 \$6732 \$7142 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1322 \$153 \$7690 \$6913 \$7608 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1323 \$16 \$6860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1324 \$16 \$7000 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1326 \$153 \$7469 \$6996 \$7142 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1327 \$16 \$7502 \$7158 \$7400 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$1328 \$16 \$7502 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1331 \$16 \$7502 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1332 \$16 \$6907 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1333 \$153 \$7336 \$6996 \$7437 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1334 \$153 \$7438 \$7236 \$6784 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1335 \$153 \$7438 \$6794 \$7437 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1336 \$153 \$7401 \$6995 \$7437 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1337 \$153 \$7402 \$6732 \$7439 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1339 \$153 \$7338 \$6794 \$7439 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1340 \$153 \$7403 \$6996 \$7439 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1341 \$153 \$7339 \$6719 \$7439 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1342 \$153 \$7471 \$7456 \$7440 \$7472 \$7470 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$1343 \$153 \$153 \$6996 \$7250 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1345 \$153 \$7340 \$7003 \$7380 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1347 \$16 \$7473 \$16 \$153 \$6909 VNB sky130_fd_sc_hd__clkbuf_2
X$1348 \$153 \$7441 \$7357 \$6797 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1349 \$153 \$7441 \$6906 \$7380 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1350 \$16 \$6754 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1351 \$16 \$6797 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1352 \$16 \$7547 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1353 \$16 \$7381 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1354 \$153 \$7457 \$7357 \$6916 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1355 \$16 \$6916 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1358 \$153 \$7457 \$6867 \$7380 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1359 \$16 \$7378 \$6990 \$7503 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$1360 \$16 \$7333 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1361 \$153 \$7383 \$7322 \$6991 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1362 \$153 \$7405 \$7322 \$6916 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1363 \$16 \$6916 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1364 \$16 \$6915 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1365 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$1367 \$153 \$7475 \$7322 \$7044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1368 \$16 \$7044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1370 \$153 \$7059 \$7323 \$6862 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1371 \$153 \$7474 \$6324 \$7382 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1372 \$153 \$7475 \$7006 \$7382 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1373 \$16 \$6797 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1376 \$153 \$7290 \$6756 \$7043 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1377 \$153 \$7406 \$6906 \$7043 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1378 \$153 \$7408 \$7476 \$7044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1379 \$16 \$7548 \$16 \$153 \$7163 VNB sky130_fd_sc_hd__clkbuf_2
X$1380 \$153 \$7504 \$7476 \$6862 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1381 \$16 \$7044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1383 \$16 \$7466 \$16 \$153 \$7458 VNB sky130_fd_sc_hd__inv_1
X$1384 \$16 \$6862 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1385 \$153 \$7409 \$6992 \$7458 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1386 \$153 \$7504 \$7003 \$7458 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1387 \$153 \$7410 \$6992 \$7316 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1388 \$153 \$7477 \$6867 \$7316 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1389 \$153 \$7478 \$7003 \$7316 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1390 \$16 \$7072 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1391 \$16 \$7212 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1392 \$16 \$6910 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1394 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$1395 \$153 \$7442 \$7479 \$6862 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1396 \$16 \$6862 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1397 \$153 \$7443 \$7384 \$6797 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1398 \$153 \$7442 \$7003 \$7612 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1399 \$153 \$7443 \$6906 \$7411 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1401 \$153 \$7480 \$6324 \$7749 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1403 \$153 \$7444 \$7384 \$6771 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1404 \$16 \$3418 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1405 \$153 \$7444 \$6865 \$7411 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1406 \$153 \$7294 \$7006 \$7411 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1408 \$153 \$7481 \$6582 \$7296 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1410 \$153 \$7752 \$7482 \$7296 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1412 \$153 \$7459 \$7327 \$7296 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1413 \$16 \$7445 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1415 \$16 \$7386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1416 \$16 \$7347 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1417 \$153 \$7483 \$6582 \$7597 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1418 \$153 \$7014 \$7484 \$7414 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$1419 \$16 \$7328 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1420 \$16 \$7484 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1422 \$16 \$7082 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1424 \$153 \$7199 \$7065 \$7257 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1425 \$16 \$7239 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1426 \$16 \$7344 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1428 \$153 \$6972 \$7551 \$7485 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$1429 \$153 \$7505 \$7550 \$7129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1431 \$16 \$7387 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1432 \$153 \$7486 \$6582 \$7388 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1434 \$153 \$7506 \$7074 \$7445 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1435 \$153 \$7506 \$7327 \$7085 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1436 \$16 \$7445 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1438 \$153 \$7086 \$8794 \$7460 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$1439 \$16 \$7495 \$7633 \$7460 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$1440 \$153 \$7487 \$7327 \$7112 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1443 \$153 \$7416 \$7366 \$7112 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1444 \$16 \$7495 \$16 \$153 \$7112 VNB sky130_fd_sc_hd__inv_1
X$1446 \$153 \$7446 \$7169 \$7328 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1447 \$153 \$7507 \$7169 \$7445 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1448 \$153 \$7446 \$7366 \$7317 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1451 \$153 \$7367 \$7215 \$7317 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1452 \$16 \$7540 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1453 \$153 \$7488 \$7490 \$6656 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1454 \$16 \$7489 \$16 \$153 \$6656 VNB sky130_fd_sc_hd__inv_1
X$1455 \$16 \$7445 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1456 \$153 \$7447 \$7171 \$7445 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1457 \$153 \$7491 \$7490 \$7264 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1458 \$16 \$7429 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1459 \$16 \$7489 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1463 \$16 \$7328 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1464 \$153 \$7448 \$7265 \$7328 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1466 \$153 \$7448 \$7366 \$7417 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1467 \$153 \$7449 \$7265 \$7387 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1468 \$153 \$7449 \$7490 \$7417 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1469 \$16 \$7498 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1471 \$16 \$7498 \$7673 \$7461 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$1472 \$153 \$7090 \$7267 \$7461 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$1473 \$153 \$7173 \$7484 \$7450 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$1475 \$153 \$7492 \$7375 \$7451 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1476 \$153 \$7418 \$7462 \$7093 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1477 \$16 \$7386 \$16 \$153 \$7451 VNB sky130_fd_sc_hd__inv_1
X$1480 \$16 \$7307 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1481 \$16 \$7049 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1482 \$153 \$7493 \$7376 \$7451 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1483 \$153 \$7419 \$7375 \$7093 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1484 \$16 \$7353 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1485 \$16 \$7464 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1486 \$153 \$7452 \$7240 \$7464 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1487 \$153 \$7452 \$7639 \$7148 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1488 \$16 \$7377 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1490 \$16 \$7709 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1493 \$16 \$7350 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1494 \$153 \$7270 \$7463 \$7148 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1495 \$16 \$7350 \$7049 \$7494 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$1496 \$153 \$7390 \$7241 \$7464 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1497 \$16 \$7464 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1498 \$16 \$7131 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1499 \$16 \$7174 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1500 \$153 \$7508 \$7643 \$7131 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1503 \$153 \$7351 \$7607 \$7097 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1504 \$16 \$7495 \$7049 \$7509 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$1505 \$153 \$7510 \$7242 \$7377 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1506 \$16 \$7377 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1507 \$16 \$7464 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1508 \$153 \$7391 \$7243 \$7464 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1509 \$16 \$7495 \$16 \$153 \$7392 VNB sky130_fd_sc_hd__inv_1
X$1511 \$16 \$7353 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1513 \$153 \$7453 \$7243 \$7353 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1514 \$153 \$7453 \$7375 \$7392 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1515 \$16 \$7464 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1516 \$153 \$7511 \$7244 \$7464 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1517 \$16 \$7489 \$16 \$153 \$6985 VNB sky130_fd_sc_hd__inv_1
X$1519 \$153 \$7275 \$7180 \$6985 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1521 \$153 \$7512 \$7244 \$7377 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1522 \$16 \$7377 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1524 \$16 \$7307 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1525 \$16 \$7353 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1526 \$153 \$7513 \$7186 \$7353 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1527 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$1528 \$16 \$7540 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1529 \$16 \$7540 \$16 \$153 \$7318 VNB sky130_fd_sc_hd__inv_1
X$1530 \$153 \$7311 \$7180 \$7318 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1532 \$16 \$7429 \$7496 \$7514 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$1534 \$153 \$7454 \$7245 \$7464 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1535 \$16 \$7429 \$16 \$153 \$7217 VNB sky130_fd_sc_hd__inv_1
X$1536 \$16 \$7307 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1537 \$16 \$6924 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1538 \$153 \$7515 \$7245 \$7307 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1539 \$153 \$5460 \$3893 \$5158 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1540 \$16 \$5158 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1542 \$16 \$7498 \$7496 \$7516 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$1544 \$153 \$7517 \$7497 \$7147 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1545 \$16 \$7498 \$16 \$153 \$7518 VNB sky130_fd_sc_hd__inv_1
X$1546 \$16 \$7498 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1547 \$16 \$4963 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1548 \$153 \$7455 \$3860 \$4963 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1549 \$153 \$5147 \$3676 \$4963 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1550 \$153 \$6964 \$5627 \$6760 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1552 \$16 \$7455 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1553 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$1554 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$1555 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$1557 \$153 \$7465 \$7544 \$7041 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1558 \$16 \$7041 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1559 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$1561 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$1563 \$153 \$7519 \$7544 \$6860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1564 \$153 \$7519 \$6732 \$7552 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1565 \$16 \$6860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1567 \$153 \$7553 \$6995 \$7552 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1568 \$16 \$7545 \$16 \$153 \$7552 VNB sky130_fd_sc_hd__inv_1
X$1569 \$153 \$7280 \$6995 \$6855 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1571 \$153 \$7499 \$6732 \$6855 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1573 \$153 \$7520 \$7053 \$6783 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1574 \$153 \$7520 \$6749 \$7137 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1575 \$16 \$7521 \$7233 \$7532 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$1576 \$153 \$7320 \$7659 \$7532 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$1577 \$16 \$7659 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1579 \$153 \$7554 \$7320 \$6981 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1580 \$16 \$7467 \$16 \$153 \$7233 VNB sky130_fd_sc_hd__clkbuf_2
X$1581 \$16 \$7521 \$16 \$153 \$7140 VNB sky130_fd_sc_hd__inv_1
X$1583 \$153 \$7555 \$7546 \$6979 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1584 \$16 \$6981 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1586 \$153 \$7501 \$6732 \$7141 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1587 \$16 \$6979 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1588 \$16 \$6860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1590 \$153 \$7248 \$6995 \$7140 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1591 \$16 \$7466 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1592 \$16 \$6733 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1593 \$153 \$7398 \$6913 \$7141 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1594 \$16 \$7466 \$7158 \$7468 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$1596 \$153 \$7533 \$7235 \$6981 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1597 \$153 \$7533 \$6930 \$7142 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1598 \$16 \$6981 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1601 \$153 \$7469 \$7235 \$7041 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1602 \$16 \$7041 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1603 \$16 \$6733 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1605 \$153 \$7522 \$7236 \$6792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1606 \$153 \$7522 \$6719 \$7437 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1607 \$153 \$7556 \$6930 \$7437 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1610 \$153 \$7557 \$7337 \$6981 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1611 \$153 \$7557 \$6930 \$7439 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1612 \$153 \$7523 \$7337 \$6783 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1613 \$153 \$7523 \$6749 \$7439 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1614 \$16 \$6783 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1615 \$16 \$7471 \$16 \$153 \$7466 VNB sky130_fd_sc_hd__clkbuf_2
X$1617 \$16 \$7558 \$16 \$153 \$7502 VNB sky130_fd_sc_hd__clkbuf_2
X$1618 \$153 \$7473 \$7472 \$7456 \$7470 \$7440 \$16 \$16 VNB
+ sky130_fd_sc_hd__nor4b_2
X$1619 \$16 \$1325 \$16 \$153 \$7559 VNB sky130_fd_sc_hd__clkbuf_2
X$1620 \$153 \$7357 \$7547 \$7591 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$1621 \$16 \$7560 \$16 \$153 \$6935 VNB sky130_fd_sc_hd__clkbuf_2
X$1622 \$16 \$1325 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1623 \$153 \$7524 \$7357 \$6754 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1625 \$153 \$7524 \$6756 \$7380 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1627 \$153 \$7525 \$7357 \$7060 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1628 \$153 \$7525 \$6324 \$7380 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1629 \$153 \$7322 \$7333 \$7503 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$1630 \$16 \$7378 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1631 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$1634 \$16 \$7378 \$16 \$153 \$7382 VNB sky130_fd_sc_hd__inv_1
X$1635 \$16 \$6991 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1636 \$16 \$7378 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1637 \$153 \$7561 \$7006 \$7562 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1638 \$153 \$7474 \$7322 \$7060 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1639 \$16 \$7548 \$16 \$153 \$6990 VNB sky130_fd_sc_hd__clkbuf_2
X$1640 \$153 \$7323 \$7659 \$7592 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$1641 \$16 \$7060 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1643 \$16 \$7521 \$16 \$153 \$7043 VNB sky130_fd_sc_hd__inv_1
X$1645 \$153 \$7563 \$7323 \$6991 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1646 \$153 \$7564 \$7323 \$6916 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1647 \$16 \$7502 \$7163 \$7407 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$1649 \$16 \$6797 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1650 \$153 \$7565 \$7476 \$6797 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1652 \$153 \$7566 \$7476 \$6916 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1653 \$153 \$7565 \$6906 \$7458 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1654 \$16 \$6916 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1655 \$16 \$7466 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1656 \$16 \$7000 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1657 \$153 \$7534 \$6324 \$7458 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1658 \$153 \$7477 \$7238 \$6916 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1660 \$16 \$6916 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1661 \$153 \$7526 \$7238 \$7060 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1662 \$153 \$7526 \$6324 \$7316 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1663 \$16 \$7060 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1664 \$16 \$7535 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1666 \$153 \$7567 \$7479 \$6797 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1667 \$16 \$6797 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1668 \$16 \$5932 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1669 \$16 \$7535 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1670 \$16 \$6753 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1673 \$16 \$6753 \$16 \$153 \$7411 VNB sky130_fd_sc_hd__inv_1
X$1674 \$153 \$7568 \$7384 \$6916 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1675 \$153 \$7569 \$7384 \$7060 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1676 \$16 \$7060 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1677 \$16 \$7342 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1678 \$153 \$7570 \$7384 \$6862 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1680 \$16 \$3418 \$7342 \$16 \$153 \$4983 VNB sky130_fd_sc_hd__and2b_2
X$1682 \$153 \$7481 \$7549 \$7067 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1683 \$153 \$7459 \$7549 \$7445 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1684 \$153 \$7385 \$7549 \$7029 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1686 \$16 \$7386 \$7633 \$7596 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$1687 \$16 \$7067 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1688 \$153 \$7483 \$7632 \$7067 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1690 \$153 \$7536 \$7482 \$7597 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1691 \$153 \$7536 \$7632 \$7239 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1692 \$16 \$7350 \$7633 \$7485 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$1693 \$16 \$7239 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1696 \$153 \$7527 \$7550 \$7239 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1697 \$153 \$7527 \$7482 \$7388 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1698 \$16 \$7445 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1699 \$153 \$7528 \$7550 \$7445 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1700 \$153 \$7528 \$7327 \$7388 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1702 \$16 \$8869 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1704 \$153 \$7074 \$8869 \$7415 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$1705 \$153 \$7487 \$7086 \$7445 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1706 \$153 \$7537 \$7215 \$7571 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1708 \$16 \$7328 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1709 \$16 \$7495 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1711 \$16 \$7445 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1712 \$153 \$7538 \$7327 \$6656 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1715 \$16 \$7387 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1716 \$153 \$7539 \$7169 \$7387 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1718 \$16 \$7540 \$7673 \$7572 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$1719 \$153 \$7488 \$7170 \$7387 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1720 \$153 \$7169 \$7693 \$7572 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$1723 \$153 \$7598 \$7171 \$7328 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1724 \$16 \$7328 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1725 \$16 \$7429 \$16 \$153 \$7264 VNB sky130_fd_sc_hd__inv_1
X$1726 \$153 \$7171 \$7614 \$7599 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$1728 \$153 \$7573 \$7265 \$7129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1730 \$16 \$7387 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1733 \$153 \$7302 \$7066 \$7417 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1735 \$16 \$7431 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1736 \$16 \$7431 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1737 \$16 \$7445 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1738 \$153 \$7529 \$7265 \$7445 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1739 \$153 \$7529 \$7327 \$7417 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1741 \$16 \$7386 \$7049 \$7574 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$1742 \$153 \$7575 \$7607 \$7451 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1745 \$153 \$7576 \$7541 \$7147 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1746 \$153 \$7576 \$7463 \$7451 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1747 \$16 \$7602 \$16 \$153 \$7489 VNB sky130_fd_sc_hd__clkbuf_2
X$1748 \$16 \$7147 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1750 \$153 \$7493 \$7541 \$7174 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1751 \$16 \$7174 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1752 \$16 \$7464 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1753 \$16 \$7353 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1756 \$16 \$8869 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1758 \$16 \$7131 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1759 \$16 \$7353 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1760 \$153 \$7420 \$7607 \$7148 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1761 \$153 \$7604 \$7240 \$7353 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1762 \$16 \$7903 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1764 \$16 \$7551 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1765 \$16 \$7049 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1766 \$153 \$7241 \$7551 \$7494 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$1768 \$16 \$7377 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1770 \$153 \$7421 \$7462 \$7148 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1772 \$153 \$7577 \$7643 \$7174 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1774 \$16 \$8794 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1775 \$16 \$7353 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1776 \$153 \$7542 \$7375 \$7149 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1777 \$153 \$7542 \$7242 \$7353 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1779 \$16 \$7464 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1780 \$16 \$7495 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1781 \$16 \$7049 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1782 \$16 \$7307 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1783 \$153 \$7578 \$7243 \$7307 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1784 \$16 \$7495 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1785 \$16 \$7377 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1786 \$153 \$7530 \$7243 \$7377 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1787 \$153 \$7530 \$7462 \$7392 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1789 \$16 \$7686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1791 \$153 \$7244 \$7686 \$7579 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$1793 \$16 \$7307 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1794 \$153 \$7543 \$7208 \$7580 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1795 \$153 \$7531 \$7688 \$7307 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1796 \$153 \$7186 \$7693 \$7426 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$1799 \$153 \$7581 \$7186 \$7464 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1800 \$153 \$7209 \$7376 \$7318 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1801 \$153 \$7245 \$7614 \$7514 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$1802 \$16 \$7431 \$7496 \$7582 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$1803 \$16 \$7267 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1804 \$153 \$6552 \$5074 \$6924 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1806 \$153 \$6369 \$5635 \$6924 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1807 \$16 \$6924 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1809 \$153 \$7187 \$7267 \$7516 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$1810 \$153 \$7583 \$7497 \$7133 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1811 \$16 \$7147 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1812 \$153 \$7277 \$7463 \$7518 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1813 \$16 \$7133 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1816 \$16 \$7498 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1817 \$16 \$7174 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1818 \$16 \$4963 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1819 \$153 \$7584 \$7497 \$7174 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1820 \$153 \$7119 \$5074 \$6760 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1821 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$1822 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$1823 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$1824 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$1825 \$153 \$9877 \$9875 \$8580 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1827 \$153 \$10056 \$8638 \$9728 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1828 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$1829 \$153 \$10030 \$10088 \$10006 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1830 \$16 \$8436 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1831 \$16 \$8114 \$16 \$153 \$9728 VNB sky130_fd_sc_hd__inv_1
X$1833 \$16 \$9026 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1834 \$16 \$8114 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1836 \$153 \$9993 \$9831 \$8580 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1838 \$153 \$9993 \$8194 \$9729 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1839 \$16 \$8580 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1840 \$16 \$8436 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1841 \$16 \$8139 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1842 \$16 \$8828 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1843 \$153 \$9603 \$9832 \$8436 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1846 \$153 \$9962 \$8912 \$9583 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1847 \$16 \$8436 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1849 \$153 \$10012 \$8638 \$9583 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1850 \$153 \$10031 \$9879 \$8580 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1851 \$16 \$8580 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1852 \$16 \$8335 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1853 \$153 \$9879 \$8335 \$9896 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$1855 \$16 \$8144 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1856 \$153 \$9963 \$8912 \$9865 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1857 \$16 \$8828 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1858 \$153 \$9994 \$9765 \$8580 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1860 \$153 \$9994 \$8194 \$9740 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1862 \$153 \$10032 \$9793 \$8580 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1864 \$153 \$9767 \$8457 \$9321 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1865 \$153 \$9964 \$8912 \$9866 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1866 \$153 \$10013 \$8737 \$9836 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1867 \$153 \$10033 \$9880 \$8828 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1868 \$153 \$9965 \$8194 \$9836 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1869 \$16 \$8715 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1870 \$16 \$8580 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1872 \$153 \$10033 \$8885 \$9836 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1873 \$153 \$10014 \$8638 \$9836 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1874 \$16 \$8828 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1875 \$16 \$8828 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1876 \$16 \$8580 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1877 \$16 \$8715 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1878 \$153 \$10034 \$9838 \$8580 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1879 \$153 \$10015 \$8638 \$9867 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1881 \$16 \$9026 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1882 \$16 \$9339 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1884 \$153 \$10034 \$8194 \$9867 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1885 \$153 \$10016 \$8726 \$9867 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1886 \$153 \$10017 \$8209 \$9867 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1888 \$153 \$10035 \$8340 \$8912 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1889 \$153 \$9770 \$8737 \$9567 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1890 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1893 \$16 \$8737 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1894 \$153 \$9968 \$8277 \$9451 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1895 \$153 \$10036 \$3696 \$9947 \$10120 \$9569 \$8957 \$10007 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$1896 \$153 \$10036 \$3306 \$9807 \$10018 \$10008 \$8806 \$10007 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$1897 \$16 \$8114 \$16 \$153 \$9868 VNB sky130_fd_sc_hd__inv_1
X$1899 \$153 \$9949 \$9900 \$8556 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1900 \$16 \$8686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1901 \$16 \$8556 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1902 \$153 \$9930 \$8727 \$9902 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1903 \$153 \$9995 \$9794 \$8686 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1904 \$153 \$9995 \$8651 \$9902 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1905 \$16 \$8686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1907 \$16 \$8886 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1908 \$16 \$8335 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1910 \$153 \$9996 \$9795 \$8686 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1911 \$153 \$9996 \$8651 \$9720 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1912 \$16 \$8686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1913 \$16 \$8503 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1914 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$1915 \$153 \$10037 \$9796 \$8686 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1916 \$16 \$8686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1918 \$153 \$10038 \$9796 \$8890 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1919 \$153 \$9812 \$9811 \$8556 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1920 \$16 \$8177 \$16 \$153 \$9586 VNB sky130_fd_sc_hd__inv_1
X$1921 \$16 \$8556 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1922 \$16 \$8177 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1924 \$153 \$10039 \$9884 \$8886 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1926 \$153 \$10019 \$8804 \$9815 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1927 \$153 \$9924 \$8651 \$9815 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1929 \$16 \$8118 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1930 \$153 \$10020 \$8789 \$9815 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1931 \$16 \$8898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1933 \$153 \$10041 \$9846 \$8686 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1934 \$16 \$8686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1935 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$1938 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$1940 \$153 \$9998 \$9846 \$8886 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1941 \$16 \$8886 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1943 \$16 \$8651 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1944 \$153 \$9997 \$8556 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$1945 \$16 \$9997 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1947 \$16 \$10042 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1948 \$16 \$10043 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1950 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1951 \$153 \$10044 \$8340 \$8610 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1952 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1953 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1954 \$153 \$9999 \$8340 \$8614 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1956 \$153 \$10040 \$8340 \$9278 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1959 \$153 \$10046 \$9732 \$8936 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1960 \$16 \$8301 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1961 \$16 \$8936 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1962 \$16 \$9275 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1963 \$16 \$9214 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1964 \$153 \$9908 \$9732 \$9214 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1965 \$153 \$9944 \$10021 \$8807 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1967 \$153 \$10021 \$8719 \$9973 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$1968 \$16 \$8673 \$16 \$153 \$10216 VNB sky130_fd_sc_hd__inv_1
X$1969 \$16 \$9214 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1971 \$16 \$8807 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1972 \$153 \$9870 \$10000 \$8807 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1973 \$153 \$10000 \$8820 \$10059 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$1974 \$16 \$8313 \$16 \$153 \$9871 VNB sky130_fd_sc_hd__inv_1
X$1977 \$153 \$9887 \$9674 \$9214 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1979 \$153 \$9888 \$9674 \$9275 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1980 \$153 \$10083 \$8627 \$10060 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$1981 \$153 \$9852 \$8842 \$9642 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1983 \$153 \$10047 \$9934 \$8936 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1984 \$153 \$10047 \$8842 \$9927 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1985 \$16 \$9642 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1987 \$16 \$8936 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1988 \$153 \$10001 \$10022 \$8936 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1989 \$153 \$10001 \$8842 \$10009 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1992 \$16 \$9045 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$1993 \$153 \$10023 \$9133 \$10009 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1994 \$153 \$10002 \$10024 \$9045 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$1995 \$153 \$10002 \$9174 \$10104 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$1997 \$16 \$8428 \$16 \$153 \$10104 VNB sky130_fd_sc_hd__inv_1
X$1998 \$153 \$9889 \$9755 \$9214 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2000 \$16 \$8666 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2002 \$153 \$9976 \$9252 \$9725 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2003 \$16 \$9188 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2004 \$153 \$10003 \$9755 \$9188 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2005 \$153 \$10003 \$8917 \$9725 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2006 \$16 \$9188 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2007 \$153 \$10010 \$8705 \$9977 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$2010 \$153 \$9892 \$9758 \$9214 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2011 \$153 \$9939 \$10010 \$8936 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2012 \$153 \$10048 \$9758 \$8807 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2013 \$16 \$8807 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2014 \$16 \$8807 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2016 \$16 \$10044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2019 \$153 \$9978 \$8842 \$9823 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2021 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2022 \$153 \$10049 \$8340 \$8923 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2023 \$153 \$10050 \$9913 \$8893 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2024 \$153 \$9980 \$8977 \$9981 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2025 \$16 \$9035 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2028 \$153 \$9893 \$9913 \$8879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2029 \$153 \$9982 \$8965 \$9981 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2030 \$16 \$8879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2031 \$153 \$10051 \$9940 \$8893 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2032 \$153 \$9914 \$8996 \$9759 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2033 \$16 \$8313 \$16 \$153 \$10108 VNB sky130_fd_sc_hd__inv_1
X$2037 \$16 \$9997 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2038 \$153 \$9985 \$8965 \$10108 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2039 \$153 \$9997 \$8893 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$2040 \$16 \$8626 \$9675 \$9986 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$2041 \$16 \$7996 \$16 \$153 \$10011 VNB sky130_fd_sc_hd__inv_1
X$2042 \$153 \$9957 \$10025 \$8893 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2044 \$153 \$10026 \$8965 \$10011 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2046 \$16 \$8626 \$16 \$153 \$10110 VNB sky130_fd_sc_hd__inv_1
X$2047 \$153 \$10052 \$10085 \$9154 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2048 \$153 \$10004 \$10085 \$8893 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2049 \$153 \$10004 \$8996 \$10110 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2050 \$16 \$9154 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2053 \$153 \$9915 \$9122 \$9708 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2054 \$153 \$10027 \$8996 \$9988 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2056 \$153 \$10053 \$10111 \$8844 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2057 \$16 \$8893 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2058 \$16 \$8844 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2059 \$153 \$9960 \$9860 \$8844 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2061 \$153 \$9918 \$9860 \$8927 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2062 \$16 \$8353 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2063 \$153 \$10028 \$8353 \$9989 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$2064 \$16 \$8879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2065 \$16 \$8844 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2066 \$153 \$10054 \$10028 \$8844 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2067 \$16 \$8666 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2071 \$16 \$8704 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2073 \$16 \$8893 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2074 \$153 \$8329 \$7463 \$8266 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2075 \$153 \$10029 \$8965 \$10005 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2076 \$153 \$8630 \$7208 \$8777 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2077 \$153 \$10055 \$9792 \$8844 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2078 \$16 \$8844 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2079 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$2081 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$2082 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$2083 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$2084 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$2085 \$16 \$8715 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2086 \$153 \$10056 \$9875 \$8715 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2089 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$2091 \$153 \$9735 \$9875 \$8436 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2092 \$153 \$10086 \$10318 \$10006 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2094 \$153 \$10057 \$9831 \$8436 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2095 \$153 \$10062 \$8885 \$9729 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2097 \$153 \$10062 \$9831 \$8828 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2098 \$153 \$9679 \$9832 \$8580 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2099 \$153 \$10087 \$10088 \$10210 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2100 \$16 \$8580 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2101 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$2102 \$153 \$10117 \$8726 \$9865 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2104 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$2105 \$153 \$10031 \$8194 \$9865 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2107 \$153 \$10089 \$9879 \$8828 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2108 \$153 \$10089 \$8885 \$9865 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2109 \$153 \$10178 \$8209 \$9865 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2110 \$16 \$8271 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2113 \$153 \$10090 \$8885 \$9740 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2114 \$16 \$8580 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2116 \$16 \$8715 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2117 \$153 \$10091 \$9793 \$8715 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2118 \$153 \$10092 \$9793 \$9026 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2119 \$153 \$10032 \$8194 \$9866 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2122 \$153 \$8838 \$8580 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$2123 \$16 \$8838 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2125 \$153 \$10014 \$9880 \$8715 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2127 \$153 \$10058 \$9838 \$8828 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2129 \$153 \$10015 \$9838 \$8715 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2130 \$16 \$8839 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2132 \$16 \$9227 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2133 \$153 \$10016 \$9838 \$9026 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2134 \$16 \$8950 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2136 \$153 \$10093 \$8340 \$8885 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2138 \$153 \$10094 \$8340 \$8194 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2139 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2140 \$153 \$10036 \$4134 \$10035 \$10079 \$10080 \$9336 \$10007 \$16 \$16
+ VNB sky130_fd_sc_hd__mux4_1
X$2141 \$16 \$8114 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2142 \$153 \$9808 \$8727 \$9451 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2143 \$16 \$7949 \$16 \$153 \$10036 VNB sky130_fd_sc_hd__clkbuf_2
X$2144 \$16 \$7949 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2146 \$16 \$7884 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2148 \$153 \$10095 \$9900 \$8647 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2149 \$153 \$9948 \$9900 \$8686 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2150 \$153 \$9882 \$9900 \$8728 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2151 \$16 \$8728 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2152 \$16 \$8728 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2155 \$153 \$10063 \$9794 \$8556 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2156 \$153 \$10063 \$8610 \$9902 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2157 \$16 \$8556 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2158 \$16 \$8271 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2159 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$2160 \$153 \$10064 \$9795 \$8886 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2162 \$16 \$8816 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2163 \$16 \$8886 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2164 \$16 \$8423 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2167 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$2168 \$153 \$10065 \$9796 \$8886 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2169 \$16 \$8886 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2170 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$2171 \$153 \$10037 \$8651 \$9842 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2172 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$2173 \$16 \$8890 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2174 \$153 \$10066 \$9811 \$8686 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2176 \$153 \$10065 \$8727 \$9842 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2177 \$16 \$8686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2178 \$16 \$8760 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2180 \$153 \$10019 \$9884 \$8816 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2181 \$16 \$8816 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2182 \$16 \$8634 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2183 \$16 \$10081 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2184 \$153 \$10020 \$9884 \$8898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2185 \$16 \$7934 \$16 \$153 \$10082 VNB sky130_fd_sc_hd__clkbuf_2
X$2187 \$16 \$7934 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2188 \$16 \$10151 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2189 \$153 \$10067 \$9846 \$8898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2190 \$153 \$10096 \$8277 \$9815 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2191 \$16 \$8898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2192 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$2193 \$153 \$10068 \$9846 \$8816 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2194 \$16 \$8816 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2195 \$16 \$10205 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2196 \$16 \$8804 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2198 \$16 \$10097 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2199 \$16 \$10098 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2200 \$16 \$10401 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2201 \$153 \$9745 \$8651 \$9746 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2202 \$153 \$10043 \$8647 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$2203 \$153 \$10069 \$8340 \$8651 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2204 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2206 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2208 \$153 \$10045 \$8340 \$8818 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2209 \$153 \$10153 \$8340 \$8676 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2211 \$153 \$8301 \$9214 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$2212 \$16 \$8818 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2216 \$16 \$9045 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2217 \$153 \$10099 \$10021 \$9045 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2218 \$16 \$8807 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2219 \$16 \$9188 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2220 \$16 \$8936 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2221 \$153 \$10100 \$10021 \$8936 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2222 \$153 \$9950 \$8917 \$9453 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2223 \$16 \$8676 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2224 \$16 \$8917 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2225 \$16 \$8936 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2227 \$153 \$10100 \$8842 \$10216 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2228 \$16 \$8313 \$9518 \$10059 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$2229 \$153 \$10102 \$10000 \$8936 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2230 \$16 \$9214 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2232 \$16 \$8807 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2233 \$153 \$9952 \$10083 \$8807 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2234 \$16 \$7996 \$9518 \$10060 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$2236 \$153 \$10070 \$10083 \$8936 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2237 \$16 \$8627 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2238 \$16 \$9031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2239 \$16 \$8936 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2240 \$153 \$9954 \$9934 \$9031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2241 \$16 \$8626 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2243 \$153 \$10103 \$9174 \$9927 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2244 \$16 \$9188 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2246 \$16 \$8807 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2248 \$153 \$10071 \$10022 \$8807 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2249 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$2250 \$16 \$9031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2251 \$16 \$8624 \$16 \$153 \$10009 VNB sky130_fd_sc_hd__inv_1
X$2252 \$153 \$10023 \$10022 \$9031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2253 \$153 \$10072 \$10024 \$8807 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2255 \$16 \$8807 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2256 \$16 \$9031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2257 \$16 \$8428 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2258 \$16 \$8936 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2259 \$153 \$10073 \$10024 \$8936 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2260 \$153 \$10073 \$8842 \$10104 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2261 \$16 \$8936 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2262 \$153 \$10105 \$10157 \$8936 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2264 \$16 \$8353 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2265 \$16 \$8165 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2268 \$16 \$9031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2270 \$16 \$8705 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2271 \$16 \$9253 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2272 \$153 \$10157 \$8353 \$9911 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$2273 \$16 \$8704 \$16 \$153 \$9872 VNB sky130_fd_sc_hd__inv_1
X$2275 \$16 \$9214 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2276 \$153 \$10106 \$8917 \$9955 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2277 \$153 \$10126 \$9174 \$9955 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2279 \$153 \$10074 \$8676 \$9955 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2281 \$153 \$10074 \$10010 \$8807 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2282 \$16 \$10045 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2283 \$16 \$9999 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2284 \$16 \$10123 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2285 \$16 \$10061 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2286 \$153 \$10075 \$4203 \$9999 \$10061 \$10084 \$9979 \$10220 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$2287 \$153 \$10048 \$8676 \$9823 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2288 \$16 \$8927 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2290 \$153 \$10107 \$9913 \$8927 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2291 \$153 \$10050 \$8996 \$9981 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2292 \$153 \$10076 \$9913 \$9034 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2293 \$153 \$10076 \$9059 \$9981 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2295 \$16 \$9154 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2296 \$16 \$9154 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2299 \$16 \$9034 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2300 \$16 \$8820 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2301 \$16 \$10043 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2302 \$153 \$10051 \$8996 \$10108 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2303 \$153 \$10043 \$8844 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$2305 \$153 \$10025 \$8627 \$9984 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$2306 \$16 \$8627 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2308 \$16 \$8626 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2310 \$16 \$8731 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2311 \$16 \$8844 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2312 \$153 \$10109 \$8977 \$10011 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2314 \$153 \$10026 \$10025 \$8844 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2315 \$16 \$8626 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2316 \$16 \$8844 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2317 \$153 \$9959 \$10085 \$8844 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2318 \$16 \$8429 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2319 \$16 \$8893 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2320 \$16 \$9035 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2322 \$153 \$10052 \$9103 \$10110 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2323 \$16 \$9134 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2325 \$153 \$10111 \$8702 \$9987 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$2326 \$153 \$10077 \$10111 \$9154 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2327 \$153 \$10077 \$9103 \$9988 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2328 \$16 \$8844 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2329 \$16 \$8927 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2332 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$2333 \$153 \$10053 \$8965 \$9988 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2334 \$16 \$9154 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2335 \$153 \$8405 \$7375 \$7076 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2336 \$153 \$10078 \$9860 \$9154 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2337 \$153 \$10078 \$9103 \$9961 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2338 \$16 \$8927 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2339 \$16 \$8704 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2341 \$16 \$9154 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2343 \$153 \$10113 \$10028 \$9154 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2344 \$153 \$10114 \$10028 \$8893 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2345 \$16 \$8704 \$16 \$153 \$10112 VNB sky130_fd_sc_hd__inv_1
X$2347 \$153 \$10115 \$9991 \$8893 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2348 \$16 \$8428 \$16 \$153 \$10005 VNB sky130_fd_sc_hd__inv_1
X$2351 \$16 \$8428 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2352 \$16 \$8844 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2353 \$16 \$9154 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2354 \$153 \$10029 \$9991 \$8844 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2355 \$153 \$8881 \$7607 \$8777 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2356 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$2357 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$2358 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$2359 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$2361 \$153 \$6049 \$5896 \$5245 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2362 \$153 \$5990 \$5174 \$5837 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2363 \$153 \$6049 \$5107 \$5837 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2364 \$153 \$6050 \$5055 \$5837 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2365 \$16 \$4320 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2366 \$16 \$6051 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2368 \$16 \$5274 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2369 \$153 \$6024 \$5896 \$5404 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2370 \$153 \$6024 \$5177 \$5837 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2371 \$16 \$5404 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2372 \$16 \$5518 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2373 \$153 \$6025 \$5976 \$5489 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2374 \$153 \$6025 \$5373 \$5977 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2376 \$153 \$5944 \$5463 \$5977 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2377 \$16 \$5489 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2378 \$16 \$6051 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2380 \$153 \$6052 \$5177 \$5977 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2381 \$153 \$6026 \$6053 \$5274 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2382 \$153 \$6054 \$5373 \$6043 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2383 \$16 \$4479 \$16 \$153 \$6043 VNB sky130_fd_sc_hd__inv_1
X$2384 \$16 \$5274 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2385 \$16 \$4616 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2388 \$153 \$6055 \$5107 \$6043 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2389 \$16 \$4896 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2390 \$16 \$5181 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2391 \$153 \$5978 \$6056 \$5181 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2392 \$153 \$6027 \$6056 \$5404 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2393 \$153 \$6027 \$5177 \$5993 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2394 \$16 \$6057 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2396 \$16 \$4421 \$16 \$153 \$5993 VNB sky130_fd_sc_hd__inv_1
X$2397 \$153 \$6028 \$5948 \$5404 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2399 \$153 \$6028 \$5177 \$6143 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2400 \$153 \$5995 \$5405 \$6143 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2401 \$16 \$4600 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2402 \$16 \$5349 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2404 \$16 \$5230 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2405 \$16 \$5245 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2406 \$153 \$6058 \$5405 \$5890 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2408 \$16 \$5181 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2409 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$2410 \$16 \$5489 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2411 \$153 \$6059 \$5874 \$5489 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2412 \$16 \$5245 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2414 \$16 \$4146 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2415 \$16 \$5518 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2416 \$153 \$6029 \$6120 \$5518 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2417 \$153 \$6029 \$5463 \$6044 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2421 \$153 \$6060 \$5065 \$6223 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$2422 \$16 \$5274 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2423 \$16 \$5245 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2424 \$153 \$6030 \$6060 \$5245 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2425 \$153 \$6030 \$5107 \$6045 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2426 \$153 \$5923 \$5373 \$5722 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2427 \$16 \$4712 \$16 \$153 \$6045 VNB sky130_fd_sc_hd__inv_1
X$2429 \$153 \$5979 \$5832 \$5518 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2430 \$153 \$5924 \$5055 \$5722 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2431 \$16 \$5518 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2432 \$153 \$6031 \$5833 \$5324 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2434 \$153 \$6031 \$5096 \$5877 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2435 \$16 \$5324 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2438 \$16 \$5467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2440 \$153 \$5997 \$5833 \$5232 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2441 \$153 \$5953 \$5287 \$5877 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2442 \$16 \$5232 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2444 \$153 \$5998 \$5901 \$5232 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2445 \$16 \$5232 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2446 \$16 \$5338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2447 \$16 \$5469 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2448 \$16 \$5080 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2450 \$153 \$6083 \$5901 \$5478 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2451 \$153 \$6061 \$5901 \$5566 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2452 \$16 \$5566 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2453 \$16 \$4479 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2454 \$153 \$6062 \$5846 \$5324 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2455 \$16 \$4479 \$16 \$153 \$6032 VNB sky130_fd_sc_hd__inv_1
X$2458 \$16 \$5478 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2459 \$16 \$5324 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2460 \$153 \$6033 \$5846 \$5271 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2461 \$153 \$6033 \$5069 \$6032 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2462 \$16 \$5271 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2463 \$153 \$6000 \$5849 \$5324 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2464 \$153 \$5957 \$5069 \$5980 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2466 \$153 \$6063 \$5849 \$5338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2467 \$153 \$6063 \$5209 \$5980 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2468 \$16 \$5338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2469 \$16 \$4146 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2470 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$2471 \$16 \$4494 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2472 \$16 \$4631 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2473 \$16 \$5109 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2474 \$153 \$5981 \$5929 \$5271 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2475 \$16 \$5271 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2477 \$16 \$4494 \$5479 \$6064 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$2478 \$153 \$6034 \$4631 \$6064 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$2479 \$153 \$6002 \$6123 \$5478 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2480 \$16 \$5478 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2482 \$16 \$4869 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2483 \$153 \$6084 \$6123 \$5324 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2485 \$16 \$4869 \$5479 \$6065 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$2486 \$153 \$6085 \$5228 \$6065 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$2488 \$153 \$6066 \$5830 \$5467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2489 \$16 \$5467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2490 \$153 \$6003 \$5390 \$5815 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2491 \$153 \$6066 \$5406 \$5815 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2493 \$153 \$6004 \$5830 \$5324 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2494 \$16 \$5271 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2495 \$16 \$5324 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2496 \$16 \$5338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2497 \$153 \$6068 \$6067 \$5819 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2499 \$153 \$6086 \$6067 \$5714 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2502 \$16 \$5819 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2503 \$16 \$5834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2504 \$153 \$6035 \$6067 \$5834 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2505 \$153 \$6035 \$5881 \$6005 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2506 \$153 \$6069 \$5470 \$6136 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2507 \$16 \$4590 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2508 \$153 \$6195 \$4590 \$6232 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$2509 \$16 \$4930 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2511 \$16 \$5856 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2512 \$16 \$5796 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2513 \$153 \$6087 \$5961 \$5796 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2515 \$153 \$6006 \$6200 \$5891 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2516 \$153 \$6087 \$5775 \$5891 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2517 \$153 \$6088 \$5961 \$5834 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2521 \$16 \$5714 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2522 \$16 \$5528 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2523 \$153 \$6036 \$5973 \$5528 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2524 \$153 \$6036 \$5500 \$6089 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2525 \$16 \$5702 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2526 \$16 \$5796 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2527 \$153 \$6037 \$5973 \$5796 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2528 \$16 \$4415 \$16 \$153 \$6089 VNB sky130_fd_sc_hd__inv_1
X$2530 \$16 \$5834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2532 \$153 \$6037 \$5775 \$6089 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2533 \$153 \$6038 \$6011 \$5834 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2534 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$2535 \$153 \$6038 \$5881 \$5985 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2536 \$153 \$6009 \$5795 \$5985 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2537 \$153 \$6010 \$5755 \$5985 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2540 \$153 \$5986 \$6011 \$5605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2542 \$16 \$5714 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2543 \$153 \$5884 \$6012 \$5714 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2544 \$16 \$5702 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2545 \$16 \$5796 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2546 \$153 \$6070 \$6012 \$5796 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2549 \$153 \$6071 \$5881 \$5892 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2550 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$2551 \$16 \$5834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2552 \$153 \$6014 \$6072 \$5834 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2553 \$153 \$6073 \$6072 \$5605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2554 \$153 \$6073 \$5625 \$5987 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2556 \$153 \$6072 \$4316 \$6015 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$2557 \$16 \$4316 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2558 \$16 \$4125 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2560 \$153 \$6016 \$5775 \$5987 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2561 \$16 \$4376 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2562 \$16 \$5718 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2563 \$153 \$6074 \$5907 \$5718 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2564 \$16 \$4954 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2565 \$16 \$4093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2566 \$16 \$4324 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2567 \$16 \$4324 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2569 \$153 \$6017 \$5575 \$5823 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2570 \$153 \$6075 \$5627 \$5823 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2572 \$16 \$5963 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2573 \$16 \$5718 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2574 \$16 \$5579 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2575 \$153 \$6039 \$6076 \$5579 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2576 \$153 \$6039 \$5484 \$6018 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2577 \$16 \$4415 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2578 \$16 \$5543 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2579 \$16 \$5887 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2581 \$153 \$6077 \$5938 \$6018 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2582 \$153 \$6046 \$5074 \$6018 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2584 \$153 \$6090 \$5717 \$5786 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2586 \$16 \$1485 \$16 \$153 \$6078 VNB sky130_fd_sc_hd__clkbuf_2
X$2588 \$153 \$6079 \$5635 \$6047 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2589 \$16 \$4415 \$5485 \$6091 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$2592 \$153 \$5866 \$5627 \$5611 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2594 \$16 \$4415 \$16 \$153 \$6048 VNB sky130_fd_sc_hd__inv_1
X$2595 \$153 \$6080 \$5635 \$6048 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2596 \$153 \$6081 \$6169 \$5609 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2597 \$16 \$5636 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2598 \$153 \$6040 \$5835 \$5636 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2601 \$153 \$6040 \$5509 \$5867 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2602 \$16 \$6078 \$16 \$153 \$5582 VNB sky130_fd_sc_hd__clkbuf_2
X$2603 \$16 \$5579 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2604 \$153 \$5912 \$5910 \$5579 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2605 \$16 \$4258 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2606 \$16 \$5609 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2607 \$153 \$6041 \$5910 \$5609 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2608 \$16 \$4464 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2611 \$153 \$6041 \$5074 \$5893 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2613 \$16 \$4464 \$16 \$153 \$5894 VNB sky130_fd_sc_hd__inv_1
X$2614 \$16 \$4464 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2615 \$153 \$6082 \$5806 \$5894 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2616 \$153 \$5914 \$5941 \$5887 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2617 \$153 \$6021 \$5484 \$5894 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2618 \$16 \$4376 \$5582 \$6022 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$2619 \$16 \$5963 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2622 \$153 \$6042 \$6023 \$5963 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2623 \$153 \$6042 \$5806 \$5895 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2624 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$2626 \$16 \$5786 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2627 \$153 \$6092 \$6023 \$5786 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2628 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$2631 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$2632 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$2633 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$2634 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$2635 \$153 \$6050 \$5896 \$5736 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2637 \$16 \$5181 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2638 \$16 \$5736 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2641 \$153 \$5917 \$5405 \$5837 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2642 \$16 \$4579 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2643 \$16 \$6051 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2644 \$153 \$5975 \$5896 \$5274 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2646 \$153 \$6093 \$5896 \$5489 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2647 \$153 \$6093 \$5373 \$5837 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2650 \$153 \$6094 \$5976 \$5274 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2651 \$153 \$6094 \$4706 \$5977 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2652 \$153 \$6095 \$5976 \$5181 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2653 \$153 \$6095 \$5174 \$5977 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2654 \$16 \$5080 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2655 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$2657 \$153 \$6055 \$6053 \$5245 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2658 \$153 \$6126 \$5174 \$6043 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2659 \$16 \$5245 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2660 \$16 \$4479 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2661 \$153 \$5919 \$5055 \$6043 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2662 \$153 \$6127 \$5463 \$5993 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2663 \$153 \$6128 \$5055 \$5993 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2665 \$16 \$4621 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2666 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$2667 \$16 \$5274 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2668 \$153 \$5994 \$6056 \$5274 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2670 \$16 \$6057 \$16 \$153 \$1433 VNB sky130_fd_sc_hd__clkbuf_2
X$2671 \$153 \$6096 \$5948 \$5274 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2672 \$153 \$6096 \$4706 \$6143 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2673 \$16 \$4600 \$16 \$153 \$6143 VNB sky130_fd_sc_hd__inv_1
X$2675 \$153 \$6144 \$5948 \$5245 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2677 \$153 \$6058 \$5874 \$5403 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2679 \$153 \$6129 \$5174 \$5890 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2680 \$16 \$5403 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2682 \$153 \$6059 \$5373 \$5890 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2685 \$153 \$6145 \$6120 \$5736 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2686 \$16 \$4869 \$5630 \$5996 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$2687 \$16 \$4869 \$16 \$153 \$6044 VNB sky130_fd_sc_hd__inv_1
X$2688 \$153 \$6097 \$6120 \$5181 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2689 \$153 \$6097 \$5174 \$6044 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2690 \$16 \$5274 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2691 \$16 \$4869 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2694 \$16 \$5065 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2695 \$16 \$5403 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2696 \$153 \$6130 \$4706 \$6045 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2697 \$153 \$6146 \$6060 \$5403 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2698 \$153 \$6098 \$6060 \$5518 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2699 \$153 \$6098 \$5463 \$6045 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2700 \$16 \$5518 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2702 \$153 \$6147 \$6121 \$5467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2703 \$153 \$5876 \$5406 \$5877 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2704 \$16 \$4742 \$16 \$153 \$6149 VNB sky130_fd_sc_hd__inv_1
X$2705 \$16 \$5324 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2706 \$153 \$6099 \$5833 \$5566 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2707 \$153 \$6099 \$5519 \$5877 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2710 \$16 \$5566 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2712 \$153 \$5968 \$5901 \$5469 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2713 \$153 \$6131 \$5287 \$6149 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2714 \$153 \$5999 \$5901 \$5467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2715 \$153 \$6083 \$5390 \$5845 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2716 \$16 \$5478 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2719 \$16 \$5467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2720 \$16 \$4896 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2721 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$2722 \$153 \$5848 \$5846 \$5467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2723 \$153 \$6061 \$5519 \$5845 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2724 \$16 \$5467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2725 \$153 \$6100 \$5846 \$5338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2726 \$16 \$5338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2727 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$2729 \$153 \$6100 \$5209 \$6032 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2730 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$2731 \$16 \$5324 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2732 \$153 \$6132 \$5390 \$5980 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2733 \$153 \$6101 \$5849 \$5467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2734 \$153 \$6101 \$5406 \$5980 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2735 \$16 \$5467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2736 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$2739 \$153 \$6102 \$5929 \$5232 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2740 \$153 \$6102 \$5205 \$5852 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2741 \$16 \$4600 \$16 \$153 \$6122 VNB sky130_fd_sc_hd__inv_1
X$2742 \$16 \$5232 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2743 \$153 \$6123 \$5109 \$6152 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$2744 \$16 \$5026 \$16 \$153 \$5982 VNB sky130_fd_sc_hd__inv_1
X$2745 \$153 \$6133 \$5287 \$5982 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2747 \$153 \$5983 \$6123 \$5271 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2748 \$153 \$5984 \$6123 \$5467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2749 \$153 \$6084 \$5096 \$5982 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2750 \$153 \$6134 \$5519 \$5982 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2751 \$16 \$5467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2752 \$16 \$4712 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2755 \$153 \$6154 \$6085 \$5467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2756 \$16 \$4869 \$16 \$153 \$6175 VNB sky130_fd_sc_hd__inv_1
X$2758 \$16 \$5469 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2759 \$153 \$6103 \$6085 \$5338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2760 \$153 \$6103 \$5209 \$6175 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2761 \$153 \$6135 \$7215 \$5932 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2763 \$153 \$6156 \$6067 \$5796 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2764 \$153 \$6068 \$6200 \$6005 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2766 \$153 \$6104 \$6195 \$5714 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2767 \$153 \$6104 \$5755 \$6136 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2768 \$16 \$5351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2770 \$16 \$5856 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2772 \$153 \$6105 \$6195 \$5856 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2773 \$153 \$6105 \$5795 \$6136 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2774 \$16 \$4780 \$16 \$153 \$6136 VNB sky130_fd_sc_hd__inv_1
X$2776 \$153 \$6106 \$5961 \$5856 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2778 \$153 \$6106 \$5795 \$5891 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2781 \$16 \$4780 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2782 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$2783 \$16 \$5714 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2784 \$153 \$6159 \$5961 \$5714 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2785 \$153 \$6088 \$5881 \$5891 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2786 \$153 \$6007 \$5973 \$5714 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2787 \$16 \$6124 \$16 \$153 \$5428 VNB sky130_fd_sc_hd__clkbuf_2
X$2789 \$16 \$4542 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2792 \$16 \$5605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2793 \$153 \$6107 \$5973 \$5605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2794 \$153 \$6107 \$5625 \$6089 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2795 \$153 \$6008 \$5470 \$6089 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2797 \$153 \$6162 \$6011 \$5819 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2798 \$16 \$4562 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2801 \$16 \$4882 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2803 \$16 \$5702 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2804 \$153 \$6164 \$6011 \$5702 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2805 \$153 \$6108 \$6011 \$5528 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2806 \$153 \$6108 \$5500 \$5985 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2807 \$153 \$6125 \$5470 \$5892 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2809 \$153 \$6125 \$6012 \$5702 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2810 \$153 \$6071 \$6012 \$5834 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2811 \$16 \$5834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2812 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$2813 \$16 \$5856 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2814 \$153 \$6109 \$6072 \$5856 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2817 \$153 \$6109 \$5795 \$5987 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2818 \$153 \$5988 \$6072 \$5702 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2819 \$16 \$5714 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2820 \$16 \$5528 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2821 \$153 \$6110 \$6072 \$5528 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2822 \$153 \$6110 \$5500 \$5987 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2825 \$16 \$4092 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2826 \$16 \$5579 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2827 \$153 \$6111 \$5907 \$5579 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2828 \$153 \$6111 \$5484 \$5823 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2829 \$16 \$4780 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2830 \$153 \$6112 \$5907 \$5963 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2831 \$153 \$6112 \$5806 \$5823 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2833 \$153 \$6077 \$6076 \$5718 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2834 \$153 \$6137 \$5806 \$6018 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2835 \$16 \$5767 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2836 \$153 \$6113 \$6076 \$5767 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2837 \$153 \$6113 \$5575 \$6018 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2838 \$16 \$5579 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2839 \$16 \$5786 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2841 \$153 \$5865 \$5484 \$5475 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2843 \$16 \$6078 \$16 \$153 \$5485 VNB sky130_fd_sc_hd__clkbuf_2
X$2844 \$153 \$6169 \$4542 \$6091 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$2845 \$153 \$6114 \$6169 \$5579 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2846 \$153 \$6114 \$5484 \$6048 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2847 \$16 \$5609 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2850 \$16 \$4542 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2851 \$16 \$4415 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2852 \$16 \$5767 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2853 \$153 \$6138 \$5509 \$6048 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2854 \$153 \$6115 \$5835 \$5767 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2855 \$153 \$6115 \$5575 \$5867 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2856 \$153 \$6116 \$5910 \$5963 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2858 \$153 \$6116 \$5806 \$5893 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2860 \$16 \$5381 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2861 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$2862 \$153 \$6020 \$5509 \$5893 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2864 \$16 \$5636 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2865 \$153 \$6117 \$5941 \$5636 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2866 \$153 \$6117 \$5509 \$5894 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2867 \$16 \$5767 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2869 \$153 \$6118 \$5941 \$5767 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2870 \$153 \$6118 \$5575 \$5894 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2872 \$16 \$5579 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2873 \$153 \$6119 \$6023 \$5579 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2874 \$153 \$6119 \$5484 \$5895 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2875 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$2877 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$2878 \$16 \$5887 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2879 \$153 \$5989 \$6023 \$5887 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2880 \$153 \$6092 \$5635 \$5895 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2881 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$2882 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$2883 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$2884 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$2886 \$153 \$7355 \$6749 \$6855 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2887 \$153 \$7919 \$6930 \$7765 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2888 \$153 \$7736 \$6930 \$7552 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2889 \$16 \$7041 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2890 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$2892 \$153 \$7794 \$6913 \$7765 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2893 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$2895 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$2896 \$153 \$7795 \$6995 \$7765 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2897 \$16 \$6979 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2899 \$153 \$7815 \$7784 \$6784 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2900 \$153 \$7712 \$7784 \$6792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2901 \$16 \$6792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2902 \$16 \$6784 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2904 \$16 \$7816 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2906 \$153 \$7796 \$6995 \$7711 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2907 \$16 \$8003 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2908 \$16 \$7816 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2909 \$153 \$7766 \$7620 \$7041 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2910 \$153 \$7766 \$6996 \$7587 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2911 \$16 \$7041 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2912 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$2913 \$16 \$7922 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2914 \$153 \$7739 \$6749 \$7587 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2917 \$153 \$7817 \$7546 \$6860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2918 \$153 \$7334 \$6732 \$7140 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2919 \$16 \$6860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2920 \$16 \$6733 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2921 \$153 \$7818 \$7546 \$6784 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2922 \$153 \$7135 \$6913 \$6733 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2923 \$16 \$6907 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2925 \$16 \$7663 \$8195 \$7819 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$2926 \$16 \$6784 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2928 \$153 \$7741 \$7701 \$6979 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2929 \$153 \$7820 \$7701 \$6860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2930 \$153 \$7767 \$7703 \$6979 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2933 \$153 \$7767 \$6995 \$7768 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2934 \$153 \$7821 \$7703 \$6784 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2935 \$153 \$7236 \$6887 \$7797 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$2937 \$16 \$7769 \$16 \$153 \$7545 VNB sky130_fd_sc_hd__clkbuf_2
X$2938 \$153 \$7798 \$7785 \$7770 \$7771 \$7705 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$2941 \$153 \$7799 \$7771 \$7770 \$7785 \$7705 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$2942 \$153 \$7771 \$7785 \$7822 \$7705 \$7770 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$2943 \$153 \$7702 \$6719 \$7772 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2944 \$16 \$7786 \$16 \$153 \$7472 VNB sky130_fd_sc_hd__clkbuf_2
X$2945 \$153 \$7456 \$7470 \$7560 \$7472 \$7440 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$2946 \$16 \$7440 \$7470 \$7456 \$7472 \$16 \$153 \$7823 VNB
+ sky130_fd_sc_hd__and4_2
X$2947 \$16 \$7288 \$16 \$153 \$7800 VNB sky130_fd_sc_hd__clkbuf_2
X$2949 \$16 \$4360 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2951 \$16 \$7656 \$16 \$153 \$7867 VNB sky130_fd_sc_hd__clkbuf_2
X$2952 \$16 \$3384 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2954 \$153 \$7610 \$7624 \$6991 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2955 \$16 \$7801 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2956 \$16 \$7656 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2958 \$153 \$7743 \$6906 \$7611 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2959 \$153 \$7657 \$7003 \$7611 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2961 \$153 \$7802 \$7006 \$7787 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2963 \$153 \$7626 \$7624 \$6916 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2964 \$16 \$6916 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2965 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$2967 \$153 \$7561 \$7627 \$7044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2968 \$153 \$7658 \$6992 \$7562 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2969 \$16 \$7044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2970 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$2972 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$2973 \$16 \$6754 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2974 \$153 \$7824 \$7707 \$6771 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2975 \$153 \$7773 \$7707 \$6991 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2976 \$153 \$7773 \$6992 \$7718 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2977 \$16 \$6991 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2979 \$16 \$7335 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2980 \$16 \$7060 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2982 \$16 \$7502 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2983 \$16 \$6797 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2984 \$153 \$7803 \$6756 \$7718 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$2985 \$153 \$7825 \$7684 \$7044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2986 \$16 \$7044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2987 \$16 \$6862 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2988 \$16 \$7466 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2989 \$16 \$8177 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2990 \$153 \$7826 \$7684 \$6754 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2991 \$16 \$6754 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$2994 \$153 \$7719 \$7788 \$7044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2995 \$153 \$7827 \$7788 \$6754 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2996 \$153 \$7774 \$7788 \$6797 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$2998 \$16 \$7663 \$16 \$153 \$7612 VNB sky130_fd_sc_hd__inv_1
X$3000 \$16 \$6754 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3004 \$16 \$7535 \$7804 \$7828 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$3005 \$153 \$7664 \$7479 \$7044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3006 \$153 \$7662 \$6867 \$7612 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3007 \$16 \$6771 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3009 \$153 \$7480 \$7708 \$7060 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3010 \$16 \$6754 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3011 \$16 \$7412 \$16 \$153 \$7829 VNB sky130_fd_sc_hd__clkbuf_2
X$3013 \$153 \$7805 \$6867 \$7749 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3014 \$16 \$6991 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3015 \$153 \$7830 \$7708 \$6991 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3016 \$153 \$7722 \$7708 \$6771 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3017 \$153 \$7751 \$7003 \$7749 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3018 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$3020 \$153 \$7775 \$7549 \$7129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3021 \$16 \$7793 \$7633 \$7776 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$3022 \$153 \$7549 \$7852 \$7776 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$3023 \$16 \$7129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3025 \$16 \$7328 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3026 \$153 \$7831 \$7632 \$7328 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3028 \$153 \$7832 \$7632 \$7129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3029 \$153 \$7632 \$7903 \$7806 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$3031 \$153 \$7724 \$7550 \$7328 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3032 \$153 \$8013 \$7215 \$7789 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3034 \$153 \$7486 \$7550 \$7067 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3035 \$16 \$7667 \$7633 \$7754 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$3036 \$16 \$7387 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3037 \$153 \$7670 \$7635 \$7239 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3038 \$16 \$7833 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3040 \$153 \$7755 \$7490 \$7571 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3041 \$16 \$8675 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3042 \$16 \$7834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3045 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$3046 \$16 \$7067 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3047 \$153 \$7637 \$7636 \$7067 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3048 \$153 \$7756 \$7490 \$7613 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3049 \$16 \$7445 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3050 \$153 \$7835 \$7636 \$7445 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3052 \$16 \$7691 \$7673 \$7836 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$3055 \$16 \$7877 \$16 \$153 \$7673 VNB sky130_fd_sc_hd__clkbuf_2
X$3056 \$16 \$7067 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3057 \$153 \$7777 \$7790 \$7067 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3059 \$153 \$7777 \$6582 \$7726 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3060 \$153 \$7727 \$7790 \$7387 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3061 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$3062 \$16 \$7029 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3064 \$16 \$7328 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3065 \$153 \$7778 \$7638 \$7328 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3067 \$153 \$7778 \$7366 \$7728 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3069 \$16 \$7695 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3070 \$153 \$7807 \$6582 \$7728 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3071 \$153 \$7808 \$7638 \$7239 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3073 \$153 \$7808 \$7482 \$7728 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3074 \$16 \$7779 \$16 \$153 \$7498 VNB sky130_fd_sc_hd__clkbuf_2
X$3075 \$153 \$7779 \$7791 \$7881 \$7792 \$7880 \$16 \$16 VNB
+ sky130_fd_sc_hd__nor4b_2
X$3077 \$16 \$7780 \$16 \$153 \$7344 VNB sky130_fd_sc_hd__clkbuf_2
X$3078 \$153 \$7837 \$7541 \$7377 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3079 \$153 \$7757 \$7180 \$7451 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3082 \$16 \$7793 \$7049 \$7838 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$3083 \$153 \$7781 \$7642 \$7147 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3084 \$153 \$7781 \$7463 \$7731 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3085 \$16 \$7464 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3086 \$153 \$7732 \$7642 \$7307 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3087 \$16 \$7307 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3088 \$16 \$7839 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3090 \$16 \$7131 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3094 \$16 \$7377 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3095 \$153 \$7643 \$7903 \$7809 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$3096 \$153 \$7733 \$7643 \$7147 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3097 \$16 \$7709 \$16 \$153 \$7734 VNB sky130_fd_sc_hd__inv_1
X$3099 \$16 \$7464 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3100 \$153 \$7840 \$7643 \$7464 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3103 \$153 \$7242 \$7668 \$7810 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$3104 \$16 \$7667 \$16 \$153 \$7149 VNB sky130_fd_sc_hd__inv_1
X$3105 \$153 \$7735 \$7242 \$7147 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3106 \$16 \$7147 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3108 \$16 \$7307 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3109 \$16 \$7147 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3110 \$153 \$7644 \$7710 \$7307 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3112 \$153 \$7811 \$7463 \$7616 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3113 \$153 \$7812 \$7710 \$7131 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3114 \$16 \$7131 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3115 \$16 \$6985 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3116 \$16 \$8291 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3117 \$16 \$7131 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3118 \$153 \$7543 \$7688 \$7131 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3119 \$16 \$7952 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3120 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$3123 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$3124 \$153 \$7813 \$7462 \$7580 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3125 \$153 \$7759 \$7180 \$7580 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3126 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$3127 \$16 \$7133 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3128 \$153 \$7841 \$7698 \$7133 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3129 \$153 \$7427 \$7462 \$7318 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3130 \$16 \$7174 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3134 \$16 \$7306 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3135 \$153 \$7231 \$7463 \$7217 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3136 \$153 \$7783 \$7208 \$7782 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3137 \$153 \$7783 \$7647 \$7131 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3138 \$16 \$7131 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3139 \$153 \$7497 \$8101 \$7814 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$3140 \$16 \$7133 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3142 \$153 \$7842 \$7647 \$7133 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3143 \$16 \$7353 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3144 \$153 \$7843 \$7497 \$7131 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3145 \$153 \$7844 \$7497 \$7377 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3146 \$16 \$7377 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3147 \$16 \$7695 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3150 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$3151 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$3152 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$3153 \$153 \$7845 \$7864 \$7041 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3154 \$153 \$7845 \$6996 \$7765 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3158 \$153 \$7883 \$7864 \$6860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3159 \$16 \$6860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3161 \$153 \$7846 \$7864 \$6792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3162 \$153 \$7846 \$6719 \$7765 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3163 \$16 \$6792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3164 \$153 \$7500 \$6913 \$7140 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3166 \$16 \$7884 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3167 \$16 \$8001 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3168 \$153 \$7815 \$6794 \$7711 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3169 \$153 \$7847 \$7784 \$6981 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3170 \$153 \$7847 \$6930 \$7711 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3171 \$153 \$7737 \$6913 \$7711 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3172 \$153 \$7865 \$6732 \$7587 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3175 \$153 \$7885 \$7620 \$6792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3176 \$16 \$6792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3177 \$16 \$7922 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3178 \$153 \$7651 \$7866 \$6860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3179 \$153 \$7886 \$7866 \$6979 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3180 \$16 \$6979 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3182 \$153 \$6863 \$6732 \$6733 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3183 \$153 \$7704 \$7866 \$6907 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3184 \$153 \$7546 \$7887 \$7819 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$3186 \$153 \$7848 \$7701 \$6783 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3188 \$153 \$7963 \$6719 \$7609 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3189 \$16 \$6783 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3190 \$16 \$6784 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3191 \$153 \$7849 \$7703 \$6981 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3193 \$153 \$7849 \$6930 \$7768 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3194 \$153 \$7742 \$6913 \$7768 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3195 \$16 \$7535 \$8195 \$7797 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$3196 \$16 \$7535 \$16 \$153 \$7437 VNB sky130_fd_sc_hd__inv_1
X$3198 \$153 \$7821 \$6794 \$7768 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3199 \$16 \$7799 \$16 \$153 \$7381 VNB sky130_fd_sc_hd__clkbuf_2
X$3200 \$16 \$7798 \$16 \$153 \$6988 VNB sky130_fd_sc_hd__clkbuf_2
X$3201 \$153 \$7769 \$7785 \$7771 \$7705 \$7770 \$16 \$16 VNB
+ sky130_fd_sc_hd__nor4b_2
X$3202 \$16 \$7945 \$6903 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$3203 \$16 \$7786 \$16 \$153 \$7785 VNB sky130_fd_sc_hd__clkbuf_2
X$3204 \$153 \$7785 \$7705 \$7888 \$7771 \$7770 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$3205 \$153 \$7741 \$6995 \$7772 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3206 \$16 \$6667 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3209 \$16 \$7889 \$16 \$153 \$7456 VNB sky130_fd_sc_hd__clkbuf_2
X$3210 \$16 \$6667 \$16 \$153 \$7786 VNB sky130_fd_sc_hd__clkbuf_2
X$3211 \$16 \$7859 \$7800 \$7867 \$153 \$7706 \$16 VNB sky130_fd_sc_hd__and3b_4
X$3212 \$153 \$7859 \$7867 \$7890 \$7800 \$16 \$16 VNB sky130_fd_sc_hd__nor3b_4
X$3213 \$16 \$7801 \$16 \$153 \$7859 VNB sky130_fd_sc_hd__clkbuf_2
X$3214 \$16 \$7823 \$16 \$153 \$7071 VNB sky130_fd_sc_hd__clkbuf_2
X$3215 \$16 \$7891 \$16 \$153 \$8037 VNB sky130_fd_sc_hd__clkbuf_2
X$3217 \$153 \$7868 \$7003 \$7787 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3219 \$16 \$5477 \$16 \$153 \$7949 VNB sky130_fd_sc_hd__clkbuf_2
X$3220 \$16 \$6451 \$16 \$153 \$7934 VNB sky130_fd_sc_hd__clkbuf_2
X$3221 \$153 \$7802 \$7946 \$7044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3223 \$153 \$7850 \$7624 \$7044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3225 \$153 \$7869 \$6324 \$7611 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3226 \$16 \$7044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3228 \$16 \$8003 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3230 \$153 \$7850 \$7006 \$7611 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3231 \$16 \$8003 \$16 \$153 \$7562 VNB sky130_fd_sc_hd__inv_1
X$3232 \$153 \$7892 \$6867 \$7562 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3234 \$153 \$7870 \$6865 \$7562 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3235 \$153 \$7745 \$6906 \$7562 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3236 \$153 \$7717 \$7707 \$6916 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3238 \$153 \$7824 \$6865 \$7718 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3239 \$153 \$7660 \$6865 \$7043 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3240 \$153 \$7803 \$7707 \$6754 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3241 \$153 \$7893 \$7707 \$7060 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3242 \$16 \$7894 \$16 \$153 \$7548 VNB sky130_fd_sc_hd__clkbuf_2
X$3243 \$16 \$7894 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3245 \$16 \$8177 \$16 \$153 \$7895 VNB sky130_fd_sc_hd__inv_1
X$3246 \$16 \$7060 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3248 \$153 \$7896 \$7684 \$6797 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3249 \$16 \$6797 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3250 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$3251 \$16 \$8118 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3252 \$153 \$7851 \$7788 \$6916 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3253 \$153 \$7851 \$6867 \$7720 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3254 \$16 \$6916 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3256 \$16 \$7887 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3257 \$153 \$7827 \$6756 \$7720 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3258 \$16 \$6771 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3259 \$16 \$6797 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3260 \$153 \$7897 \$7479 \$6771 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3262 \$153 \$7384 \$6903 \$7899 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$3263 \$153 \$7898 \$7006 \$8260 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3266 \$153 \$7871 \$7708 \$6754 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3267 \$153 \$7805 \$7708 \$6916 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3268 \$153 \$7871 \$6756 \$7749 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3269 \$16 \$7288 \$16 \$153 \$7872 VNB sky130_fd_sc_hd__clkbuf_2
X$3270 \$16 \$6862 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3271 \$153 \$7295 \$7490 \$5932 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3273 \$153 \$7830 \$6992 \$7749 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3275 \$16 \$7387 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3276 \$153 \$7900 \$7549 \$7387 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3277 \$16 \$5932 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3278 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$3280 \$153 \$7873 \$7065 \$7860 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3281 \$153 \$7901 \$7215 \$7860 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3282 \$16 \$7793 \$16 \$153 \$7296 VNB sky130_fd_sc_hd__inv_1
X$3284 \$16 \$7852 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3285 \$16 \$7129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3286 \$153 \$7902 \$7874 \$7129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3287 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$3288 \$16 \$7709 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3289 \$16 \$7129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3290 \$153 \$7831 \$7366 \$7597 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3291 \$16 \$7445 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3292 \$16 \$7709 \$7633 \$7806 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$3294 \$153 \$7875 \$7065 \$7924 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3295 \$16 \$7903 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3297 \$16 \$7387 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3298 \$153 \$7723 \$7550 \$7387 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3299 \$153 \$7861 \$6582 \$7789 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3300 \$153 \$7853 \$7876 \$7082 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3301 \$153 \$7853 \$7065 \$7789 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3302 \$16 \$7239 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3303 \$16 \$7667 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3305 \$16 \$7877 \$16 \$153 \$7633 VNB sky130_fd_sc_hd__clkbuf_2
X$3306 \$16 \$7445 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3307 \$153 \$7878 \$6582 \$7571 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3308 \$153 \$7905 \$7635 \$7445 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3309 \$16 \$7904 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3310 \$16 \$7328 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3311 \$153 \$7906 \$7636 \$7328 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3312 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$3313 \$16 \$7239 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3315 \$153 \$7907 \$7636 \$7239 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3317 \$153 \$7835 \$7327 \$7613 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3318 \$153 \$7692 \$7065 \$7613 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3319 \$153 \$7725 \$7790 \$7029 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3320 \$16 \$7029 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3322 \$16 \$7239 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3325 \$16 \$7387 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3327 \$153 \$7854 \$7790 \$7239 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3328 \$153 \$7854 \$7482 \$7726 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3330 \$153 \$7855 \$7638 \$7029 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3332 \$153 \$7855 \$7066 \$7728 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3334 \$16 \$8101 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3335 \$16 \$7067 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3336 \$153 \$7807 \$7638 \$7067 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3337 \$153 \$7638 \$8101 \$7600 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$3338 \$16 \$7879 \$16 \$153 \$7431 VNB sky130_fd_sc_hd__clkbuf_2
X$3339 \$153 \$7879 \$7791 \$7880 \$7881 \$7792 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$3340 \$16 \$7880 \$7792 \$7881 \$7791 \$16 \$153 \$7602 VNB
+ sky130_fd_sc_hd__and4_2
X$3343 \$153 \$7603 \$7208 \$7451 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3344 \$153 \$7837 \$7462 \$7451 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3345 \$153 \$7642 \$7852 \$7838 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$3346 \$16 \$7908 \$16 \$153 \$7350 VNB sky130_fd_sc_hd__clkbuf_2
X$3347 \$16 \$7793 \$16 \$153 \$7731 VNB sky130_fd_sc_hd__inv_1
X$3348 \$153 \$7910 \$7642 \$7377 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3350 \$16 \$7909 \$16 \$153 \$7793 VNB sky130_fd_sc_hd__clkbuf_2
X$3351 \$153 \$7911 \$7642 \$7353 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3352 \$16 \$7353 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3353 \$16 \$7377 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3354 \$16 \$7307 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3355 \$153 \$7677 \$7376 \$7731 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3356 \$16 \$7709 \$7049 \$7809 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$3357 \$153 \$7856 \$7643 \$7307 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3360 \$153 \$7856 \$7607 \$7734 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3361 \$153 \$7912 \$7643 \$7353 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3362 \$153 \$7840 \$7639 \$7734 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3363 \$16 \$7667 \$7049 \$7810 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$3364 \$153 \$7913 \$7862 \$7131 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3366 \$16 \$7377 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3367 \$153 \$7758 \$7607 \$7149 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3368 \$153 \$7811 \$7710 \$7147 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3369 \$153 \$7857 \$7710 \$7377 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3370 \$153 \$7857 \$7462 \$7616 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3371 \$16 \$8772 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3372 \$16 \$7353 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3375 \$16 \$7615 \$16 \$153 \$7496 VNB sky130_fd_sc_hd__clkbuf_2
X$3376 \$153 \$7914 \$7688 \$7353 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3378 \$16 \$7952 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3379 \$16 \$7174 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3380 \$153 \$7858 \$7688 \$7174 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3381 \$153 \$7858 \$7376 \$7580 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3382 \$16 \$7353 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3383 \$16 \$7915 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3387 \$16 \$7691 \$16 \$153 \$7882 VNB sky130_fd_sc_hd__inv_1
X$3388 \$16 \$7691 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3389 \$16 \$7377 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3390 \$153 \$7760 \$7463 \$7882 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3391 \$153 \$7916 \$7698 \$7377 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3392 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$3394 \$16 \$7131 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3395 \$153 \$8198 \$7863 \$7131 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3398 \$153 \$7689 \$7639 \$7782 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3399 \$153 \$7761 \$7376 \$7782 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3400 \$153 \$7917 \$7647 \$7353 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3401 \$153 \$7918 \$7647 \$7307 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3402 \$16 \$7307 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3403 \$16 \$7131 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3407 \$153 \$7210 \$7208 \$7518 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3408 \$153 \$7314 \$7462 \$7518 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3409 \$153 \$7433 \$7639 \$7518 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3410 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$3411 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$3412 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$3413 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$3414 \$153 \$2686 \$2510 \$1658 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3415 \$153 \$2687 \$2643 \$1658 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3416 \$153 \$2582 \$1792 \$2343 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3417 \$153 \$2532 \$2064 \$2343 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3419 \$16 \$1658 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3420 \$16 \$1037 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3421 \$16 \$945 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3422 \$153 \$2510 \$945 \$2668 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$3423 \$16 \$2932 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3424 \$153 \$2619 \$2377 \$1980 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3425 \$153 \$2669 \$2252 \$2110 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3426 \$153 \$2670 \$1815 \$2110 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3428 \$153 \$2433 \$2511 \$1980 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3429 \$153 \$2644 \$2252 \$2179 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3430 \$153 \$2619 \$2009 \$2179 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3431 \$153 \$2645 \$1943 \$2275 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3432 \$153 \$2584 \$2252 \$2275 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3433 \$16 \$1522 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3434 \$16 \$972 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3436 \$153 \$2621 \$2380 \$1980 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3437 \$16 \$1795 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3438 \$153 \$2646 \$1211 \$2534 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$3439 \$16 \$1980 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3440 \$16 \$1553 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3441 \$16 \$1348 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3442 \$16 \$1211 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3443 \$153 \$2688 \$2646 \$2180 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3445 \$153 \$2587 \$2646 \$1980 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3446 \$16 \$1067 \$16 \$153 \$2586 VNB sky130_fd_sc_hd__inv_1
X$3447 \$153 \$2588 \$2290 \$2024 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3448 \$153 \$2575 \$1943 \$1594 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3449 \$153 \$2621 \$2009 \$1594 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3450 \$16 \$691 \$16 \$153 \$2671 VNB sky130_fd_sc_hd__inv_1
X$3452 \$16 \$691 \$2647 \$2690 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$3454 \$153 \$2691 \$2649 \$1942 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3455 \$16 \$1942 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3456 \$16 \$2024 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3457 \$153 \$2692 \$2478 \$2024 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3458 \$16 \$1048 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3459 \$16 \$1048 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3460 \$153 \$2589 \$1792 \$2386 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3463 \$153 \$2673 \$2252 \$2741 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3464 \$153 \$2648 \$2064 \$2671 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3465 \$16 \$1658 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3467 \$153 \$2649 \$1173 \$2590 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$3468 \$153 \$2537 \$2009 \$2386 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3469 \$153 \$2672 \$2210 \$2634 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3470 \$16 \$2414 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3473 \$153 \$3120 \$1547 \$2634 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3474 \$16 \$2538 \$2650 \$2635 \$2674 \$16 \$153 \$2675 VNB
+ sky130_fd_sc_hd__and4_2
X$3475 \$16 \$2435 \$2420 \$2436 \$2434 \$16 \$153 \$2514 VNB
+ sky130_fd_sc_hd__and4_2
X$3476 \$16 \$2113 \$16 \$153 \$2635 VNB sky130_fd_sc_hd__clkbuf_2
X$3477 \$153 \$2622 \$2652 \$1923 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3479 \$153 \$2622 \$1895 \$2636 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3482 \$153 \$2651 \$1806 \$2636 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3484 \$16 \$2089 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3485 \$16 \$1923 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3486 \$16 \$585 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3487 \$16 \$2743 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3489 \$153 \$2676 \$2652 \$2043 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3490 \$153 \$2623 \$2652 \$1805 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3491 \$16 \$1348 \$2539 \$2677 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$3493 \$153 \$2678 \$1703 \$2594 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3494 \$153 \$2595 \$1954 \$2299 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3495 \$153 \$2624 \$2708 \$2042 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3496 \$16 \$2042 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3497 \$16 \$1966 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3498 \$153 \$2653 \$2555 \$2043 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3499 \$16 \$2043 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3501 \$153 \$2625 \$2555 \$1845 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3502 \$153 \$2558 \$1924 \$2557 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3503 \$16 \$2042 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3505 \$153 \$2679 \$2359 \$2089 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3506 \$16 \$2089 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3508 \$153 \$2559 \$1471 \$2499 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3510 \$153 \$2626 \$2525 \$2042 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3511 \$153 \$2680 \$1806 \$2499 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3512 \$153 \$2626 \$1924 \$2499 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3513 \$16 \$2199 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3515 \$153 \$2682 \$2597 \$2042 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3516 \$16 \$691 \$16 \$153 \$2346 VNB sky130_fd_sc_hd__inv_1
X$3518 \$153 \$2681 \$2026 \$2346 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3519 \$153 \$2682 \$1924 \$2346 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3520 \$153 \$2598 \$2200 \$1845 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3521 \$16 \$1845 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3522 \$153 \$2654 \$2026 \$2637 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3523 \$16 \$2089 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3524 \$153 \$2655 \$1924 \$2637 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3526 \$153 \$2638 \$2560 \$1923 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3527 \$153 \$2638 \$1895 \$2637 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3528 \$16 \$2199 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3529 \$16 \$1923 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3530 \$16 \$588 \$16 \$153 \$2500 VNB sky130_fd_sc_hd__inv_1
X$3531 \$153 \$2516 \$2578 \$1805 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3532 \$16 \$2042 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3533 \$16 \$1805 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3534 \$16 \$1923 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3535 \$16 \$2043 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3537 \$153 \$2693 \$2578 \$2043 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3538 \$153 \$2600 \$2026 \$2500 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3539 \$153 \$2694 \$2517 \$2016 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3540 \$153 \$2656 \$1558 \$2639 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3541 \$16 \$2016 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3542 \$16 \$902 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3543 \$16 \$1044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3545 \$153 \$2601 \$1993 \$2161 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3546 \$153 \$2602 \$1868 \$2161 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3547 \$16 \$902 \$1968 \$2603 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$3548 \$16 \$1878 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3550 \$153 \$2640 \$2485 \$1878 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3552 \$153 \$2640 \$1868 \$2502 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3553 \$16 \$1489 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3554 \$16 \$1044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3556 \$16 \$1879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3557 \$16 \$1969 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3558 \$153 \$2695 \$2485 \$1969 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3559 \$153 \$2562 \$1558 \$2502 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3560 \$16 \$1650 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3562 \$153 \$2696 \$1245 \$2657 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$3564 \$153 \$2658 \$1558 \$2641 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3566 \$16 \$1879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3567 \$16 \$1969 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3568 \$153 \$2697 \$1558 \$2627 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3569 \$16 \$2232 \$16 \$153 \$2627 VNB sky130_fd_sc_hd__inv_1
X$3570 \$16 \$2659 \$16 \$153 \$1929 VNB sky130_fd_sc_hd__clkbuf_2
X$3571 \$153 \$2604 \$2092 \$2280 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3573 \$153 \$2628 \$2309 \$2098 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3575 \$153 \$2628 \$1993 \$2334 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3577 \$153 \$2717 \$2438 \$2641 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3578 \$153 \$2683 \$1715 \$2641 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3580 \$153 \$2605 \$2579 \$2098 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3581 \$16 \$2098 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3583 \$16 \$2016 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3584 \$153 \$2607 \$2579 \$2016 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3586 \$16 \$2104 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3587 \$153 \$2565 \$2579 \$2104 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3588 \$153 \$2579 \$1719 \$2608 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$3589 \$16 \$1184 \$16 \$153 \$2606 VNB sky130_fd_sc_hd__inv_1
X$3590 \$16 \$1719 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3591 \$16 \$1184 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3592 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$3593 \$153 \$2609 \$1712 \$2188 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3596 \$16 \$2098 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3597 \$153 \$2660 \$2092 \$2504 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3598 \$16 \$1878 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3599 \$153 \$2698 \$2732 \$1878 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3600 \$153 \$2368 \$723 \$2545 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$3601 \$16 \$1120 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3603 \$16 \$2204 \$16 \$153 \$2684 VNB sky130_fd_sc_hd__clkbuf_2
X$3604 \$16 \$2793 \$16 \$153 \$2204 VNB sky130_fd_sc_hd__clkbuf_2
X$3605 \$16 \$2793 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3607 \$16 \$2576 \$16 \$153 \$2126 VNB sky130_fd_sc_hd__clkbuf_2
X$3609 \$153 \$2505 \$2337 \$2464 \$2372 \$2371 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$3610 \$16 \$2576 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3612 \$153 \$2371 \$2337 \$2611 \$2372 \$2464 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$3613 \$153 \$2699 \$2685 \$2700 \$2684 \$2733 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$3614 \$16 \$1972 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3615 \$153 \$2661 \$2056 \$2613 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3616 \$153 \$2466 \$1936 \$2402 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3618 \$153 \$2701 \$2612 \$2093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3619 \$16 \$2093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3621 \$153 \$2702 \$2612 \$1960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3622 \$16 \$1960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3624 \$16 \$2085 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3625 \$153 \$2529 \$1935 \$2085 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3628 \$16 \$1973 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3629 \$16 \$1860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3630 \$16 \$1960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3631 \$153 \$2629 \$1935 \$1960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3632 \$153 \$2629 \$2086 \$2506 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3633 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$3635 \$16 \$1860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3636 \$153 \$2507 \$2581 \$1860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3639 \$16 \$2192 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3641 \$16 \$1973 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3642 \$153 \$2630 \$2581 \$1973 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3643 \$153 \$2630 \$2056 \$2491 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3645 \$153 \$2570 \$1719 \$2550 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$3646 \$153 \$2662 \$2269 \$2508 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3650 \$153 \$2631 \$2570 \$1973 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3651 \$153 \$2631 \$2056 \$2508 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3652 \$16 \$1973 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3653 \$16 \$2085 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3654 \$153 \$2632 \$2403 \$2085 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3655 \$153 \$2615 \$2269 \$2282 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3658 \$153 \$2703 \$2403 \$2093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3659 \$153 \$2663 \$2265 \$2032 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3660 \$153 \$2663 \$2524 \$2093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3662 \$153 \$2664 \$2265 \$2178 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3663 \$16 \$508 \$16 \$153 \$2178 VNB sky130_fd_sc_hd__inv_1
X$3664 \$16 \$508 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3666 \$16 \$724 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3667 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$3668 \$153 \$2665 \$2267 \$2178 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3669 \$153 \$2666 \$2086 \$2178 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3670 \$153 \$2667 \$2056 \$2642 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3671 \$153 \$2133 \$2572 \$2031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3672 \$16 \$2031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3673 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$3676 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$3677 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$3678 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$3679 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$3680 \$153 \$2735 \$2510 \$1980 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3682 \$16 \$1658 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3683 \$16 \$1980 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3686 \$153 \$2736 \$2643 \$1942 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3687 \$153 \$2737 \$2643 \$2180 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3688 \$16 \$2180 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3690 \$16 \$1037 \$2932 \$2668 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$3691 \$153 \$2497 \$2377 \$1942 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3693 \$16 \$1942 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3695 \$16 \$1980 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3696 \$153 \$2644 \$2377 \$2180 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3697 \$16 \$2180 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3698 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$3699 \$153 \$2738 \$2511 \$2024 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3700 \$153 \$2727 \$2009 \$2886 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3701 \$16 \$2024 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3703 \$16 \$2006 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3705 \$153 \$2645 \$2511 \$2006 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3706 \$16 \$1795 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3707 \$153 \$2633 \$2380 \$2024 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3708 \$153 \$2728 \$2009 \$3149 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3709 \$153 \$2738 \$2210 \$2275 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3710 \$16 \$2024 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3711 \$16 \$2006 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3713 \$153 \$2739 \$2646 \$2006 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3714 \$16 \$1067 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3715 \$16 \$1658 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3716 \$16 \$899 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3717 \$16 \$2180 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3718 \$153 \$2740 \$2704 \$1980 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3719 \$153 \$2705 \$2704 \$1658 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3721 \$16 \$1658 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3722 \$16 \$1980 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3723 \$16 \$1980 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3724 \$16 \$2024 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3725 \$153 \$2689 \$2704 \$1795 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3726 \$153 \$2704 \$842 \$2690 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$3727 \$153 \$2706 \$1815 \$2741 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3728 \$153 \$2691 \$2064 \$2741 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3730 \$16 \$1594 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3731 \$16 \$2647 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3732 \$153 \$2692 \$2210 \$2386 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3733 \$153 \$2673 \$2649 \$2180 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3734 \$16 \$2180 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3735 \$16 \$1173 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3736 \$16 \$2647 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3737 \$16 \$1658 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3738 \$153 \$2707 \$2649 \$1658 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3739 \$16 \$1048 \$16 \$153 \$2741 VNB sky130_fd_sc_hd__inv_1
X$3741 \$153 \$2707 \$1547 \$2741 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3742 \$153 \$2742 \$1943 \$2634 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3743 \$153 \$2445 \$2674 \$2538 \$2635 \$2650 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$3744 \$153 \$2729 \$2674 \$2635 \$2650 \$2538 \$16 \$16 VNB
+ sky130_fd_sc_hd__nor4b_2
X$3745 \$16 \$2539 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3746 \$153 \$2652 \$945 \$2592 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$3748 \$16 \$2539 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3750 \$153 \$2651 \$2652 \$1965 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3751 \$16 \$1037 \$16 \$153 \$2636 VNB sky130_fd_sc_hd__inv_1
X$3752 \$153 \$2744 \$2652 \$2089 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3753 \$153 \$2745 \$2652 \$2042 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3754 \$16 \$2042 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3757 \$16 \$2043 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3758 \$153 \$2676 \$1954 \$2636 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3759 \$153 \$2708 \$1553 \$2677 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$3760 \$153 \$2709 \$2708 \$2089 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3761 \$153 \$2709 \$2026 \$2746 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3762 \$16 \$1013 \$1966 \$2554 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$3764 \$153 \$2730 \$1954 \$2746 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3765 \$153 \$2710 \$2555 \$2199 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3766 \$153 \$2556 \$2026 \$2557 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3767 \$153 \$2653 \$1954 \$2557 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3768 \$153 \$2710 \$2184 \$2557 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3769 \$16 \$2362 \$16 \$153 \$2539 VNB sky130_fd_sc_hd__clkbuf_2
X$3771 \$153 \$2747 \$2359 \$2043 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3772 \$153 \$2679 \$2026 \$2327 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3773 \$153 \$2680 \$2525 \$1965 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3774 \$153 \$2748 \$1954 \$2499 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3775 \$16 \$1965 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3776 \$16 \$2042 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3777 \$16 \$691 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3780 \$16 \$691 \$2347 \$2596 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$3781 \$153 \$2681 \$2597 \$2089 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3782 \$16 \$2089 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3783 \$16 \$2042 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3785 \$153 \$2711 \$2597 \$1805 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3786 \$153 \$2711 \$1703 \$2346 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3787 \$16 \$1805 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3788 \$16 \$1048 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3790 \$153 \$2654 \$2560 \$2089 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3791 \$16 \$1048 \$16 \$153 \$2637 VNB sky130_fd_sc_hd__inv_1
X$3792 \$153 \$2749 \$2560 \$1965 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3793 \$16 \$1965 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3794 \$153 \$2578 \$757 \$2712 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$3795 \$16 \$588 \$2347 \$2712 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$3797 \$153 \$2713 \$2578 \$2042 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3798 \$153 \$2713 \$1924 \$2500 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3799 \$153 \$2599 \$1895 \$2500 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3801 \$153 \$2693 \$1954 \$2500 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3802 \$153 \$2714 \$1471 \$2500 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3803 \$16 \$2104 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3805 \$153 \$2715 \$2517 \$2104 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3806 \$153 \$2750 \$1715 \$2639 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3807 \$153 \$2715 \$2092 \$2161 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3808 \$153 \$2773 \$2438 \$2161 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3809 \$153 \$2694 \$1715 \$2161 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3810 \$16 \$1878 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3811 \$16 \$2098 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3813 \$153 \$2751 \$2485 \$2098 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3814 \$16 \$1378 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3816 \$16 \$1879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3817 \$153 \$2716 \$2731 \$1879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3818 \$153 \$2716 \$1558 \$2752 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3819 \$153 \$2695 \$1613 \$2502 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3822 \$16 \$2016 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3823 \$153 \$2753 \$1715 \$2752 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3824 \$16 \$2232 \$1929 \$2657 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$3826 \$153 \$2697 \$2696 \$1879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3827 \$153 \$2788 \$2696 \$1969 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3828 \$16 \$2659 \$16 \$153 \$1968 VNB sky130_fd_sc_hd__clkbuf_2
X$3830 \$16 \$2105 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3833 \$153 \$2717 \$2796 \$2105 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3834 \$16 \$1929 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3835 \$16 \$901 \$1929 \$2718 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$3836 \$153 \$2796 \$998 \$2718 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$3837 \$16 \$1878 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3838 \$153 \$2719 \$2579 \$1878 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3840 \$16 \$998 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3841 \$153 \$2719 \$1868 \$2606 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3843 \$16 \$2105 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3844 \$153 \$2720 \$2579 \$2105 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3845 \$153 \$2720 \$2438 \$2606 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3846 \$153 \$2721 \$2579 \$1756 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3848 \$153 \$2721 \$1712 \$2606 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3850 \$16 \$2104 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3851 \$153 \$2660 \$2732 \$2104 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3852 \$153 \$2722 \$2732 \$2098 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3853 \$153 \$2722 \$1993 \$2504 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3854 \$16 \$1756 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3857 \$153 \$2698 \$1868 \$2504 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3858 \$153 \$2776 \$1715 \$2504 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3860 \$16 \$2936 \$16 \$153 \$2189 VNB sky130_fd_sc_hd__clkbuf_2
X$3861 \$16 \$2936 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3863 \$153 \$2519 \$2685 \$2733 \$2699 \$2684 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$3864 \$16 \$2126 \$16 \$153 \$2699 VNB sky130_fd_sc_hd__clkbuf_2
X$3865 \$16 \$1120 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3867 \$153 \$2699 \$2684 \$2723 \$2685 \$2733 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$3868 \$16 \$2754 \$16 \$153 \$1599 VNB sky130_fd_sc_hd__clkbuf_2
X$3870 \$16 \$2734 \$16 \$153 \$815 VNB sky130_fd_sc_hd__clkbuf_2
X$3871 \$16 \$2723 \$16 \$153 \$1758 VNB sky130_fd_sc_hd__clkbuf_2
X$3872 \$153 \$2755 \$2612 \$2191 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3873 \$16 \$2700 \$16 \$153 \$1514 VNB sky130_fd_sc_hd__clkbuf_2
X$3874 \$153 \$2661 \$2612 \$1973 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3875 \$153 \$2755 \$2267 \$2613 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3876 \$16 \$1973 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3879 \$153 \$2701 \$2265 \$2613 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3881 \$16 \$2232 \$1885 \$2756 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$3882 \$153 \$2757 \$2831 \$1860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3884 \$153 \$2614 \$1935 \$1973 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3885 \$16 \$901 \$1885 \$2779 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$3886 \$16 \$1885 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3890 \$16 \$901 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3891 \$16 \$901 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3893 \$153 \$2724 \$2581 \$2192 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3894 \$153 \$2724 \$2269 \$2491 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3895 \$16 \$2191 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3896 \$153 \$2758 \$2581 \$2191 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3897 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$3901 \$16 \$1960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3902 \$153 \$2725 \$2570 \$1960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3903 \$153 \$2725 \$2086 \$2508 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3905 \$16 \$2191 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3906 \$153 \$2726 \$2570 \$2191 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3907 \$153 \$2726 \$2267 \$2508 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3910 \$153 \$2804 \$700 \$2783 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$3911 \$16 \$815 \$16 \$153 \$2759 VNB sky130_fd_sc_hd__inv_1
X$3912 \$153 \$2760 \$2269 \$2759 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3913 \$16 \$2093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3914 \$153 \$2703 \$2265 \$2282 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3915 \$153 \$2761 \$1936 \$2759 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3916 \$153 \$2762 \$2271 \$2178 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3918 \$153 \$2664 \$2572 \$2093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3919 \$16 \$2093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3921 \$16 \$2191 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3922 \$153 \$2665 \$2572 \$2191 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3924 \$16 \$1973 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3925 \$153 \$2242 \$2572 \$1973 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3928 \$16 \$1960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3929 \$153 \$2666 \$2572 \$1960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3930 \$153 \$2844 \$2086 \$2642 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3931 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$3933 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$3934 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$3935 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$3936 \$153 \$5514 \$5486 \$5403 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3937 \$16 \$5403 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3938 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$3939 \$153 \$5515 \$5266 \$5518 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3941 \$153 \$5438 \$5373 \$5120 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3943 \$16 \$5518 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3945 \$16 \$3692 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3946 \$16 \$5151 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3947 \$153 \$5487 \$5200 \$5489 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3948 \$153 \$5487 \$5373 \$5166 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3950 \$153 \$5412 \$5200 \$5403 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3951 \$16 \$5403 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3952 \$16 \$3638 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3954 \$16 \$3841 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3956 \$16 \$3841 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3958 \$153 \$5516 \$5240 \$5404 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3959 \$16 \$5404 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3960 \$16 \$5518 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3962 \$16 \$3778 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3963 \$153 \$5440 \$5240 \$5489 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3964 \$153 \$5440 \$5373 \$5276 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3965 \$16 \$5489 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3966 \$16 \$5403 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3969 \$153 \$5413 \$5267 \$5489 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3970 \$16 \$5489 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3971 \$16 \$5403 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3973 \$16 \$3714 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3974 \$153 \$5441 \$5267 \$5404 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3975 \$153 \$5441 \$5177 \$5277 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3976 \$16 \$5404 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3977 \$16 \$5183 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3978 \$16 \$3714 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3979 \$16 \$5176 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3981 \$153 \$5488 \$5347 \$5404 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3982 \$16 \$5404 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3983 \$16 \$5125 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3984 \$153 \$5415 \$5347 \$5489 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3985 \$16 \$5489 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3986 \$16 \$4107 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3987 \$153 \$5416 \$5246 \$5403 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3990 \$153 \$5490 \$5373 \$5337 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3991 \$153 \$5417 \$5246 \$5404 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3992 \$16 \$5404 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3993 \$153 \$5418 \$5461 \$5274 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$3994 \$153 \$5462 \$5463 \$5337 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$3995 \$16 \$3907 \$16 \$153 \$5517 VNB sky130_fd_sc_hd__inv_1
X$3997 \$16 \$4246 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$3998 \$16 \$3886 \$5630 \$5491 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$3999 \$153 \$5466 \$4246 \$5491 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$4000 \$16 \$5518 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4001 \$153 \$5465 \$5055 \$5464 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4002 \$153 \$153 \$5405 \$5203 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4003 \$153 \$153 \$5463 \$5203 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4005 \$16 \$5463 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4006 \$16 \$3886 \$16 \$153 \$5464 VNB sky130_fd_sc_hd__inv_1
X$4008 \$153 \$5465 \$5466 \$5736 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4009 \$16 \$5736 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4011 \$16 \$5186 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4012 \$16 \$5477 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4014 \$153 \$5362 \$5128 \$5467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4015 \$153 \$5520 \$3660 \$5492 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$4016 \$16 \$5467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4018 \$153 \$5419 \$5128 \$5469 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4019 \$16 \$5478 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4021 \$153 \$5444 \$5248 \$5469 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4022 \$153 \$5444 \$5287 \$5270 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4023 \$153 \$5493 \$5519 \$5270 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4024 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$4026 \$153 \$5421 \$5248 \$5467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4027 \$16 \$5467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4029 \$16 \$5186 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4031 \$16 \$3767 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4032 \$153 \$5521 \$5350 \$5478 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4033 \$153 \$5468 \$5350 \$5469 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4035 \$16 \$5478 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4036 \$16 \$5469 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4038 \$153 \$5423 \$5253 \$5478 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4039 \$16 \$5478 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4041 \$153 \$5522 \$5253 \$5469 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4042 \$16 \$5469 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4043 \$16 \$5183 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4044 \$16 \$5186 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4045 \$153 \$5494 \$5406 \$5283 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4047 \$153 \$5523 \$5231 \$5478 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4048 \$153 \$5424 \$5231 \$5469 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4049 \$16 \$3997 \$5713 \$5524 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$4050 \$16 \$5469 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4052 \$153 \$5495 \$5254 \$5467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4054 \$16 \$3997 \$16 \$153 \$5171 VNB sky130_fd_sc_hd__inv_1
X$4055 \$16 \$5478 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4056 \$16 \$5467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4057 \$153 \$5525 \$5254 \$5469 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4058 \$16 \$3886 \$5479 \$5446 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$4059 \$16 \$5469 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4061 \$153 \$5526 \$5273 \$5469 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4062 \$153 \$5378 \$5209 \$5286 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4064 \$16 \$3907 \$5479 \$5447 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$4065 \$153 \$5392 \$5273 \$5467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4066 \$16 \$5338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4067 \$16 \$5478 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4068 \$153 \$5527 \$5407 \$5478 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4069 \$16 \$3907 \$16 \$153 \$5339 VNB sky130_fd_sc_hd__inv_1
X$4070 \$16 \$3907 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4072 \$153 \$5448 \$5205 \$5339 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4074 \$153 \$5393 \$5407 \$5338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4075 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4076 \$16 \$5338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4077 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4078 \$153 \$3278 \$1482 \$5625 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4079 \$153 \$3417 \$1482 \$5470 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4080 \$16 \$1436 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4083 \$153 \$1436 \$5528 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$4084 \$16 \$5351 \$4881 \$5449 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$4085 \$153 \$5496 \$5470 \$5471 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4086 \$16 \$4834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4087 \$153 \$5039 \$5480 \$5450 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$4088 \$16 \$4093 \$5428 \$5529 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$4090 \$153 \$5530 \$5039 \$3889 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4091 \$16 \$4093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4092 \$153 \$5041 \$5543 \$5451 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$4093 \$153 \$5427 \$5041 \$4048 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4094 \$16 \$5543 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4095 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$4097 \$153 \$5395 \$3962 \$5016 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4098 \$153 \$5497 \$5470 \$5571 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4099 \$153 \$5042 \$5379 \$5453 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$4100 \$153 \$4931 \$5498 \$5430 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$4102 \$153 \$5499 \$5500 \$5472 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4104 \$16 \$3960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4106 \$153 \$5396 \$3716 \$4992 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4107 \$153 \$4952 \$5473 \$5501 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$4108 \$153 \$5454 \$4952 \$3960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4109 \$153 \$5454 \$3716 \$5138 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4111 \$16 \$3960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4112 \$16 \$4048 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4114 \$153 \$5431 \$4920 \$4048 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4115 \$16 \$5400 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4116 \$153 \$5481 \$3716 \$4953 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4117 \$16 \$4016 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4118 \$16 \$4048 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4119 \$153 \$5432 \$5043 \$4048 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4120 \$153 \$5456 \$3716 \$5139 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4122 \$153 \$5408 \$5043 \$3889 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4124 \$153 \$4920 \$5306 \$5409 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$4126 \$16 \$5482 \$4542 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$4127 \$16 \$5482 \$4590 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$4128 \$16 \$5482 \$4047 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$4129 \$16 \$5482 \$4560 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$4130 \$16 \$5482 \$4430 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$4131 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4132 \$16 \$5435 \$16 \$153 \$5194 VNB sky130_fd_sc_hd__clkbuf_2
X$4133 \$16 \$5355 \$4784 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$4136 \$16 \$5483 \$5498 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$4137 \$16 \$5435 \$16 \$153 \$5483 VNB sky130_fd_sc_hd__clkbuf_2
X$4138 \$16 \$5483 \$4756 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$4139 \$16 \$5483 \$5480 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$4140 \$16 \$5483 \$5452 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$4142 \$153 \$3357 \$1482 \$5484 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4144 \$16 \$4760 \$5116 \$5299 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$4145 \$153 \$3273 \$1482 \$5509 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4147 \$153 \$5576 \$4276 \$5502 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$4148 \$153 \$5503 \$5074 \$5474 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4149 \$153 \$5197 \$5541 \$5504 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$4151 \$16 \$3602 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4152 \$153 \$5505 \$5484 \$5474 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4153 \$16 \$3870 \$5485 \$5531 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$4154 \$16 \$3691 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4156 \$153 \$5506 \$5074 \$5475 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4157 \$153 \$5382 \$3893 \$5019 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4159 \$153 \$5369 \$3142 \$5019 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4160 \$153 \$5533 \$4047 \$5507 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$4161 \$153 \$5198 \$5379 \$5476 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$4163 \$16 \$5331 \$5116 \$5476 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$4165 \$16 \$3898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4166 \$153 \$5370 \$5303 \$3898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4167 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$4168 \$16 \$4129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4169 \$153 \$5304 \$5198 \$4129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4171 \$153 \$5508 \$5509 \$5614 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4174 \$153 \$5163 \$5799 \$5458 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$4175 \$16 \$3826 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4176 \$153 \$5410 \$5163 \$3826 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4177 \$16 \$3567 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4178 \$16 \$5400 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4179 \$16 \$3567 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4180 \$153 \$4738 \$3986 \$3567 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4181 \$153 \$5510 \$4414 \$5011 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4183 \$153 \$5144 \$5473 \$5384 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$4184 \$16 \$4016 \$16 \$153 \$5511 VNB sky130_fd_sc_hd__inv_1
X$4185 \$153 \$4839 \$3719 \$5011 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4186 \$153 \$5534 \$5144 \$3898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4187 \$153 \$5560 \$5002 \$5512 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$4189 \$16 \$5579 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4190 \$153 \$5307 \$5199 \$3691 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4191 \$16 \$3834 \$16 \$153 \$5309 VNB sky130_fd_sc_hd__inv_1
X$4193 \$153 \$5513 \$5806 \$5309 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4194 \$16 \$3826 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4195 \$16 \$5609 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4196 \$153 \$5310 \$5560 \$5609 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4197 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$4200 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$4201 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$4202 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$4203 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$4204 \$153 \$5535 \$5486 \$5245 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4205 \$16 \$5181 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4206 \$16 \$5245 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4208 \$153 \$5437 \$5405 \$5120 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4209 \$153 \$5536 \$5486 \$5489 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4210 \$16 \$5489 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4211 \$16 \$5274 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4212 \$153 \$5439 \$5177 \$5120 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4213 \$16 \$4579 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4214 \$153 \$5486 \$3660 \$5584 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$4215 \$16 \$5489 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4217 \$16 \$3638 \$16 \$153 \$4579 VNB sky130_fd_sc_hd__inv_1
X$4218 \$153 \$5178 \$5200 \$5518 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4219 \$16 \$5518 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4221 \$153 \$5546 \$5463 \$5276 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4222 \$153 \$5546 \$5240 \$5518 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4223 \$153 \$5516 \$5177 \$5276 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4225 \$153 \$5537 \$5240 \$5403 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4226 \$153 \$5537 \$5405 \$5276 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4227 \$153 \$5414 \$5267 \$5403 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4228 \$153 \$5641 \$5201 \$5561 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$4231 \$153 \$5538 \$5267 \$5518 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4232 \$153 \$5538 \$5463 \$5277 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4233 \$16 \$5518 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4234 \$16 \$3761 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4236 \$153 \$5711 \$5125 \$5562 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$4237 \$153 \$5488 \$5177 \$5168 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4238 \$16 \$5274 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4241 \$153 \$5246 \$4107 \$5585 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$4242 \$153 \$5490 \$5246 \$5489 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4243 \$16 \$5489 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4244 \$16 \$5403 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4246 \$16 \$3658 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4247 \$153 \$5462 \$5246 \$5518 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4248 \$16 \$5518 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4250 \$16 \$5518 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4251 \$16 \$3949 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4252 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$4253 \$153 \$5587 \$5461 \$5245 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4254 \$153 \$5588 \$5461 \$5518 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4255 \$16 \$8554 \$153 \$1482 \$16 VNB sky130_fd_sc_hd__clkbuf_4
X$4256 \$16 \$8554 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4257 \$153 \$5547 \$5177 \$5464 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4259 \$153 \$5547 \$5466 \$5404 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4260 \$16 \$5404 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4262 \$153 \$5589 \$5466 \$5518 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4263 \$153 \$5563 \$5107 \$5464 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4264 \$16 \$5518 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4266 \$153 \$5565 \$5519 \$5564 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4268 \$153 \$5590 \$5548 \$5467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4269 \$16 \$3638 \$5186 \$5492 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$4270 \$16 \$5324 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4271 \$153 \$5591 \$5548 \$5566 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4272 \$153 \$5318 \$5519 \$5169 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4273 \$16 \$5478 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4274 \$16 \$5469 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4276 \$16 \$3638 \$16 \$153 \$5564 VNB sky130_fd_sc_hd__inv_1
X$4278 \$153 \$5493 \$5248 \$5566 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4279 \$16 \$5566 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4280 \$153 \$5420 \$5248 \$5478 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4281 \$153 \$5592 \$5520 \$5232 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4282 \$16 \$5232 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4283 \$16 \$5478 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4284 \$16 \$3841 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4286 \$153 \$5593 \$5350 \$5467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4287 \$153 \$5743 \$5350 \$5566 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4288 \$16 \$5566 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4289 \$153 \$5422 \$5253 \$5467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4290 \$16 \$5467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4291 \$16 \$3761 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4292 \$16 \$3879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4295 \$153 \$5594 \$5253 \$5566 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4296 \$16 \$5566 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4298 \$16 \$4106 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4299 \$153 \$5494 \$5231 \$5467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4300 \$153 \$5523 \$5390 \$5283 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4301 \$16 \$4106 \$5713 \$5597 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$4302 \$16 \$5478 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4305 \$153 \$5254 \$4107 \$5524 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$4307 \$153 \$5425 \$5254 \$5478 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4308 \$153 \$5426 \$5254 \$5566 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4309 \$153 \$5525 \$5287 \$5171 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4311 \$16 \$5566 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4312 \$153 \$5599 \$5273 \$5566 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4313 \$153 \$5526 \$5287 \$5286 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4314 \$16 \$5469 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4316 \$153 \$5539 \$5549 \$5338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4317 \$153 \$5567 \$5096 \$5631 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4320 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$4322 \$153 \$5527 \$5390 \$5339 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4323 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$4324 \$16 \$5469 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4325 \$153 \$5540 \$5407 \$5469 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4326 \$153 \$5540 \$5287 \$5339 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4327 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$4330 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4331 \$153 \$3352 \$1482 \$6200 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4332 \$16 \$6200 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4334 \$16 \$5470 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4335 \$16 \$16 \$153 VNB sky130_fd_sc_hd__conb_1
X$4336 \$153 \$153 \$5625 \$5568 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4337 \$153 \$153 \$5470 \$5568 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4338 \$153 \$153 \$6200 \$5568 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4339 \$16 \$5351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4341 \$16 \$5541 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4342 \$153 \$5632 \$4276 \$5529 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$4343 \$16 \$4276 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4344 \$16 \$5351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4345 \$153 \$5569 \$5500 \$5340 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4346 \$16 \$3889 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4347 \$16 \$5480 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4348 \$153 \$5679 \$4196 \$5601 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$4349 \$153 \$5530 \$3962 \$5015 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4351 \$153 \$5367 \$5041 \$3960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4352 \$153 \$5570 \$5755 \$5571 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4353 \$16 \$3960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4355 \$153 \$5655 \$4126 \$5429 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$4356 \$153 \$5572 \$5500 \$5571 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4357 \$16 \$3929 \$5428 \$5551 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$4359 \$153 \$5552 \$4047 \$5551 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$4360 \$16 \$4048 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4361 \$153 \$5542 \$4931 \$3889 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4363 \$153 \$5542 \$3962 \$4992 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4365 \$16 \$5017 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4366 \$16 \$3960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4367 \$153 \$5553 \$5500 \$5624 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4369 \$16 \$4011 \$5906 \$5554 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$4370 \$153 \$5633 \$4168 \$5554 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$4371 \$153 \$5573 \$5470 \$5624 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4372 \$16 \$5702 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4373 \$153 \$5481 \$4920 \$3960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4374 \$153 \$5455 \$3962 \$4953 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4377 \$153 \$5656 \$4152 \$5604 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$4378 \$153 \$5555 \$5500 \$5727 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4380 \$16 \$3889 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4381 \$153 \$5657 \$5625 \$5434 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4382 \$153 \$5043 \$5799 \$5398 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$4383 \$16 \$3814 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4384 \$16 \$3834 \$5906 \$5556 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$4386 \$153 \$5658 \$5002 \$5556 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$4387 \$16 \$5482 \$4126 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$4388 \$16 \$5605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4389 \$153 \$5606 \$5470 \$5574 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4390 \$153 \$5634 \$4125 \$5607 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$4391 \$16 \$5483 \$5543 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$4392 \$16 \$5483 \$4759 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$4393 \$16 \$5483 \$5541 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$4394 \$16 \$5194 \$4781 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$4395 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4397 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4398 \$16 \$4957 \$16 \$153 \$5353 VNB sky130_fd_sc_hd__clkbuf_2
X$4399 \$16 \$4938 \$16 \$153 \$4882 VNB sky130_fd_sc_hd__clkbuf_2
X$4400 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4401 \$153 \$3358 \$1482 \$5575 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4402 \$16 \$4093 \$5485 \$5502 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$4404 \$153 \$5503 \$5576 \$5609 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4405 \$16 \$5351 \$5116 \$5504 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$4408 \$153 \$5505 \$5576 \$5579 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4409 \$16 \$5579 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4410 \$16 \$4139 \$5485 \$5557 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$4411 \$153 \$5532 \$4126 \$5557 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$4412 \$153 \$5610 \$5532 \$5579 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4413 \$16 \$4139 \$16 \$153 \$5611 VNB sky130_fd_sc_hd__inv_1
X$4415 \$16 \$5543 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4416 \$16 \$5379 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4417 \$16 \$5609 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4418 \$153 \$5612 \$5532 \$5609 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4419 \$153 \$5457 \$3860 \$5019 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4421 \$16 \$5963 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4422 \$153 \$5613 \$5533 \$5963 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4423 \$16 \$3929 \$16 \$153 \$5614 VNB sky130_fd_sc_hd__inv_1
X$4424 \$16 \$3929 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4428 \$16 \$5636 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4429 \$153 \$5508 \$5533 \$5636 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4430 \$16 \$4168 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4431 \$16 \$4011 \$5582 \$5558 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$4432 \$153 \$5578 \$4168 \$5558 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$4433 \$16 \$4011 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4434 \$16 \$4011 \$16 \$153 \$5559 VNB sky130_fd_sc_hd__inv_1
X$4435 \$16 \$5579 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4436 \$153 \$5577 \$5806 \$5559 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4438 \$153 \$5615 \$5578 \$5579 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4439 \$153 \$5580 \$5074 \$5559 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4440 \$16 \$5579 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4441 \$153 \$5544 \$5637 \$5579 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4442 \$153 \$5544 \$5484 \$5511 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4443 \$16 \$3898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4444 \$16 \$5609 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4446 \$153 \$5581 \$5509 \$5511 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4447 \$153 \$5617 \$4125 \$5616 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$4448 \$16 \$3834 \$5582 \$5512 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$4450 \$153 \$5545 \$5560 \$5579 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4451 \$153 \$5545 \$5484 \$5309 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4452 \$16 \$4125 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4454 \$16 \$4092 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4455 \$16 \$3834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4456 \$16 \$5636 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4457 \$153 \$5311 \$5560 \$5636 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4458 \$153 \$5583 \$5627 \$5692 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4459 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$4460 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$4461 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$4462 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$4463 \$153 \$1975 \$1873 \$2006 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4464 \$16 \$2006 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4466 \$153 \$2007 \$1873 \$1942 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4467 \$153 \$2007 \$2064 \$1762 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4468 \$16 \$1942 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4470 \$16 \$264 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4472 \$16 \$710 \$16 \$153 \$1669 VNB sky130_fd_sc_hd__inv_1
X$4473 \$16 \$531 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4475 \$16 \$2006 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4476 \$153 \$1787 \$1774 \$2006 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4477 \$153 \$2323 \$2252 \$1669 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4479 \$16 \$1595 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4481 \$16 \$1795 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4483 \$153 \$2065 \$1763 \$1980 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4485 \$153 \$2033 \$2252 \$1789 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4486 \$16 \$1980 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4488 \$153 \$2008 \$1888 \$2024 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4489 \$153 \$1889 \$1888 \$1658 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4490 \$153 \$2008 \$2210 \$1861 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4491 \$16 \$1658 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4495 \$16 \$454 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4496 \$153 \$2034 \$1943 \$1793 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4498 \$153 \$2066 \$1963 \$1980 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4499 \$153 \$2035 \$2064 \$1793 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4500 \$16 \$2006 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4501 \$153 \$2023 \$1766 \$2006 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4503 \$153 \$2023 \$1943 \$1767 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4504 \$16 \$1980 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4505 \$16 \$1942 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4506 \$16 \$2006 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4507 \$153 \$2067 \$1675 \$2006 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4508 \$153 \$1979 \$2009 \$1767 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4509 \$153 \$2036 \$1676 \$1980 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4511 \$153 \$2010 \$1676 \$1942 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4512 \$153 \$2010 \$2064 \$1670 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4514 \$16 \$2024 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4515 \$153 \$2037 \$1797 \$2024 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4516 \$153 \$2036 \$2009 \$1670 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4518 \$16 \$1508 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4520 \$153 \$2068 \$1797 \$1980 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4521 \$153 \$2037 \$2210 \$1671 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4522 \$16 \$1980 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4524 \$16 \$2025 \$16 \$153 \$264 VNB sky130_fd_sc_hd__clkbuf_2
X$4525 \$153 \$2025 \$1768 \$1777 \$1816 \$1799 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$4526 \$153 \$1816 \$1768 \$2069 \$1799 \$1777 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$4527 \$16 \$2100 \$16 \$153 \$1768 VNB sky130_fd_sc_hd__clkbuf_2
X$4530 \$16 \$377 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4531 \$153 \$2011 \$1863 \$1842 \$1875 \$2038 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$4533 \$16 \$1842 \$2038 \$1875 \$1863 \$16 \$153 \$2070 VNB
+ sky130_fd_sc_hd__and4_2
X$4534 \$16 \$2011 \$16 \$153 \$582 VNB sky130_fd_sc_hd__clkbuf_2
X$4536 \$16 \$264 \$1292 \$1982 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$4537 \$153 \$2012 \$2039 \$1923 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4538 \$153 \$2012 \$1895 \$1944 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4540 \$153 \$2071 \$1919 \$2089 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4541 \$16 \$2089 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4542 \$16 \$1923 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4543 \$153 \$1984 \$2039 \$1845 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4544 \$153 \$2072 \$1919 \$2043 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4545 \$16 \$2043 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4548 \$16 \$754 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4550 \$16 \$2089 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4552 \$16 \$541 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4553 \$153 \$2073 \$1779 \$2043 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4554 \$16 \$2043 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4555 \$16 \$2199 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4556 \$16 \$1966 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4557 \$153 \$2013 \$1921 \$1805 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4559 \$153 \$2040 \$1954 \$1922 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4561 \$153 \$2041 \$2026 \$1922 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4563 \$16 \$1923 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4564 \$153 \$2014 \$1697 \$2042 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4565 \$153 \$1985 \$1806 \$1866 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4566 \$153 \$2014 \$1924 \$1866 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4567 \$16 \$1525 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4569 \$16 \$323 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4570 \$16 \$2089 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4571 \$16 \$1965 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4574 \$16 \$535 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4575 \$16 \$356 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4577 \$16 \$842 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4578 \$153 \$1867 \$1700 \$2042 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4579 \$16 \$2042 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4580 \$16 \$356 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4582 \$153 \$2027 \$1700 \$2043 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4583 \$153 \$2027 \$1954 \$1822 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4584 \$16 \$2043 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4587 \$153 \$1986 \$1770 \$2043 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4588 \$16 \$2043 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4589 \$16 \$380 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4590 \$153 \$2074 \$1770 \$2042 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4591 \$153 \$1987 \$1780 \$2043 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4592 \$16 \$2043 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4593 \$16 \$2042 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4595 \$153 \$2015 \$1780 \$2199 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4596 \$153 \$2015 \$2184 \$1704 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4597 \$153 \$2044 \$1967 \$1923 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4598 \$153 \$1988 \$1703 \$2028 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4599 \$16 \$1805 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4600 \$16 \$1923 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4601 \$16 \$1845 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4603 \$153 \$2044 \$1895 \$2028 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4604 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4605 \$153 \$2075 \$1482 \$353 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4606 \$153 \$2076 \$1876 \$2016 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4607 \$153 \$2045 \$2092 \$1540 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4608 \$16 \$2016 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4609 \$16 \$1929 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4612 \$16 \$426 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4613 \$16 \$426 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4614 \$153 \$1955 \$1868 \$1540 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4615 \$16 \$426 \$16 \$153 \$1540 VNB sky130_fd_sc_hd__inv_1
X$4617 \$153 \$2017 \$1781 \$2105 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4618 \$153 \$2046 \$2092 \$1679 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4619 \$153 \$2017 \$2438 \$1679 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4621 \$16 \$2098 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4624 \$153 \$2077 \$1781 \$2016 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4625 \$153 \$2047 \$1993 \$1679 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4626 \$16 \$964 \$16 \$153 \$2078 VNB sky130_fd_sc_hd__inv_1
X$4627 \$153 \$2079 \$1900 \$2105 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4628 \$153 \$2048 \$2092 \$1771 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4629 \$16 \$424 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4632 \$153 \$2079 \$2438 \$1771 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4633 \$153 \$2049 \$1715 \$1771 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4634 \$16 \$1756 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4635 \$16 \$2016 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4636 \$153 \$2080 \$1880 \$2016 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4637 \$16 \$856 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4638 \$16 \$265 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4640 \$153 \$2050 \$2438 \$1674 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4642 \$16 \$798 \$16 \$153 \$1674 VNB sky130_fd_sc_hd__inv_1
X$4644 \$16 \$1969 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4645 \$153 \$1991 \$1558 \$1674 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4647 \$16 \$1878 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4648 \$153 \$1710 \$1928 \$1878 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4649 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$4650 \$16 \$1969 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4651 \$153 \$1772 \$1928 \$1969 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4653 \$16 \$151 \$16 \$153 \$1542 VNB sky130_fd_sc_hd__inv_1
X$4656 \$16 \$151 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4657 \$16 \$1627 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4658 \$16 \$306 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4659 \$16 \$2016 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4660 \$153 \$2081 \$1903 \$2016 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4661 \$16 \$1456 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4662 \$16 \$306 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4663 \$153 \$2051 \$1993 \$1759 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4664 \$153 \$1994 \$1868 \$1759 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4665 \$153 \$2052 \$2438 \$1759 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4668 \$16 \$1599 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4670 \$153 \$2018 \$2092 \$1996 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4671 \$153 \$1995 \$1613 \$1996 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4672 \$153 \$1445 \$112 \$1811 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4674 \$16 \$2053 \$16 \$153 \$80 VNB sky130_fd_sc_hd__clkbuf_2
X$4675 \$16 \$2054 \$16 \$153 \$399 VNB sky130_fd_sc_hd__clkbuf_2
X$4676 \$153 \$1882 \$1970 \$1812 \$1782 \$1831 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$4678 \$16 \$2055 \$16 \$153 \$1812 VNB sky130_fd_sc_hd__clkbuf_2
X$4679 \$16 \$1475 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4681 \$16 \$1811 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4683 \$16 \$2029 \$16 \$153 \$438 VNB sky130_fd_sc_hd__clkbuf_2
X$4684 \$153 \$2029 \$1905 \$1855 \$1883 \$1971 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$4685 \$153 \$1883 \$1905 \$2030 \$1971 \$1855 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$4686 \$16 \$2030 \$16 \$153 \$798 VNB sky130_fd_sc_hd__clkbuf_2
X$4687 \$16 \$1972 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4688 \$16 \$1811 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4689 \$16 \$1319 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4690 \$16 \$426 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4691 \$16 \$387 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4692 \$153 \$2082 \$1906 \$2031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4695 \$16 \$1973 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4696 \$153 \$1974 \$884 \$1856 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$4697 \$153 \$1998 \$2056 \$1999 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4698 \$16 \$884 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4699 \$16 \$1960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4700 \$16 \$1885 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4701 \$153 \$2083 \$1974 \$1960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4702 \$16 \$1960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4703 \$16 \$1860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4704 \$16 \$423 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4705 \$16 \$1973 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4707 \$153 \$2084 \$1974 \$1973 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4709 \$153 \$1910 \$1909 \$1960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4710 \$153 \$2057 \$2265 \$1870 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4711 \$153 \$2099 \$856 \$2019 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$4713 \$153 \$1912 \$2058 \$1973 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4714 \$16 \$1973 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4715 \$16 \$2085 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4717 \$16 \$2031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4718 \$153 \$1871 \$2058 \$2031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4719 \$153 \$2001 \$2086 \$2172 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4720 \$16 \$1973 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4722 \$16 \$829 \$1885 \$2059 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$4724 \$153 \$2004 \$948 \$2059 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$4725 \$16 \$151 \$16 \$153 \$2020 VNB sky130_fd_sc_hd__inv_1
X$4727 \$153 \$2002 \$2086 \$2020 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4728 \$16 \$2031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4729 \$16 \$2031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4730 \$153 \$2003 \$2000 \$2020 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4731 \$153 \$2021 \$2004 \$2031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4733 \$153 \$2021 \$1936 \$1940 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4734 \$153 \$2060 \$2269 \$1940 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4736 \$153 \$2005 \$2004 \$1960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4737 \$16 \$2085 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4738 \$153 \$2272 \$1938 \$2085 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4739 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$4741 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$4743 \$16 \$1973 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4744 \$153 \$2022 \$1938 \$1973 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4745 \$153 \$2061 \$2267 \$1872 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4746 \$153 \$2062 \$2269 \$1872 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4747 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$4748 \$153 \$2063 \$1936 \$2032 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4750 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$4751 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$4752 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$4753 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$4754 \$153 \$1887 \$1873 \$1980 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4755 \$16 \$1980 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4756 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$4758 \$153 \$2109 \$2009 \$2110 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4759 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$4761 \$153 \$2135 \$1873 \$2180 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4762 \$153 \$2135 \$2252 \$1762 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4763 \$153 \$2134 \$2210 \$1762 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4765 \$16 \$2024 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4767 \$16 \$279 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4769 \$153 \$2096 \$1943 \$1669 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4770 \$16 \$582 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4771 \$153 \$2033 \$1763 \$2180 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4772 \$153 \$2111 \$1815 \$1669 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4773 \$16 \$2180 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4774 \$16 \$662 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4775 \$153 \$2137 \$1888 \$1980 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4777 \$153 \$2065 \$2009 \$1789 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4778 \$16 \$2024 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4779 \$16 \$1980 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4780 \$16 \$2006 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4781 \$153 \$2034 \$1963 \$2006 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4782 \$153 \$2138 \$1963 \$2024 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4783 \$153 \$2097 \$2252 \$1793 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4785 \$16 \$2024 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4786 \$16 \$1980 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4788 \$16 \$323 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4789 \$153 \$2087 \$1766 \$2180 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4790 \$153 \$2139 \$1766 \$1942 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4792 \$153 \$2140 \$1675 \$1942 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4794 \$153 \$2112 \$1675 \$2024 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4795 \$153 \$2112 \$2210 \$1796 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4797 \$153 \$2142 \$1676 \$2024 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4799 \$153 \$2142 \$2210 \$1670 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4800 \$16 \$849 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4801 \$16 \$1659 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4803 \$16 \$1795 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4804 \$153 \$2143 \$1797 \$1942 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4805 \$16 \$1942 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4806 \$16 \$716 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4807 \$16 \$716 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4808 \$153 \$2144 \$1797 \$2180 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4809 \$153 \$2144 \$2252 \$1671 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4810 \$16 \$2180 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4812 \$16 \$685 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4813 \$16 \$585 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4815 \$16 \$1658 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4817 \$153 \$2145 \$1816 \$1777 \$1768 \$1799 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$4819 \$16 \$2113 \$16 \$153 \$1816 VNB sky130_fd_sc_hd__clkbuf_2
X$4820 \$16 \$2195 \$16 \$153 \$1799 VNB sky130_fd_sc_hd__clkbuf_2
X$4821 \$16 \$2114 \$16 \$153 \$1777 VNB sky130_fd_sc_hd__clkbuf_2
X$4822 \$16 \$2100 \$16 \$153 \$1863 VNB sky130_fd_sc_hd__clkbuf_2
X$4823 \$153 \$1981 \$2038 \$1842 \$1875 \$1863 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$4824 \$153 \$1863 \$2038 \$2101 \$1875 \$1842 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$4825 \$16 \$2101 \$16 \$153 \$1067 VNB sky130_fd_sc_hd__clkbuf_2
X$4827 \$16 \$1292 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4829 \$16 \$2115 \$16 \$153 \$899 VNB sky130_fd_sc_hd__clkbuf_2
X$4830 \$16 \$1292 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4831 \$16 \$1292 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4833 \$16 \$2199 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4834 \$16 \$1965 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4835 \$153 \$2088 \$1919 \$2199 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4836 \$153 \$1983 \$1919 \$2042 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4837 \$153 \$2071 \$2026 \$1864 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4838 \$16 \$2042 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4840 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$4841 \$153 \$2116 \$1703 \$1944 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4842 \$16 \$1845 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4843 \$153 \$2148 \$1779 \$2089 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4844 \$153 \$2149 \$1779 \$2199 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4845 \$153 \$2073 \$1954 \$1483 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4847 \$16 \$582 \$1966 \$2150 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$4849 \$153 \$2040 \$1921 \$2043 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4850 \$16 \$2043 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4851 \$16 \$1965 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4852 \$16 \$1805 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4853 \$153 \$2117 \$1697 \$2043 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4854 \$153 \$2117 \$1954 \$1866 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4855 \$16 \$2043 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4858 \$153 \$2118 \$2026 \$1866 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4860 \$16 \$849 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4861 \$16 \$1292 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4863 \$16 \$1292 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4864 \$153 \$2151 \$1820 \$2043 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4865 \$153 \$2151 \$1954 \$1844 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4866 \$153 \$2102 \$2184 \$1844 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4867 \$16 \$2043 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4868 \$16 \$849 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4870 \$153 \$2154 \$1700 \$2089 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4871 \$153 \$2154 \$2026 \$1822 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4872 \$16 \$2089 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4874 \$153 \$2155 \$1770 \$2089 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4875 \$153 \$2155 \$2026 \$1752 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4876 \$16 \$2089 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4879 \$153 \$2090 \$1770 \$2199 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4880 \$153 \$2090 \$2184 \$1752 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4881 \$16 \$2199 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4882 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$4883 \$153 \$2156 \$1780 \$2089 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4884 \$153 \$2156 \$2026 \$1704 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4886 \$153 \$2119 \$1895 \$2120 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4887 \$16 \$652 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4888 \$153 \$2121 \$2184 \$2028 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4889 \$16 \$2089 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4890 \$153 \$2157 \$1967 \$1845 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4892 \$153 \$1990 \$1806 \$2028 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4893 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$4894 \$16 \$353 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4895 \$16 \$2104 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4897 \$153 \$2045 \$1876 \$2104 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4899 \$16 \$1543 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4900 \$16 \$2105 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4901 \$16 \$2098 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4902 \$153 \$2160 \$1876 \$2098 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4903 \$153 \$2160 \$1993 \$1540 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4904 \$16 \$2104 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4905 \$16 \$387 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4907 \$16 \$2016 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4909 \$153 \$2122 \$1613 \$2161 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4911 \$153 \$2162 \$2103 \$1878 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4912 \$153 \$2047 \$1781 \$2098 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4913 \$153 \$2103 \$884 \$1946 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$4915 \$153 \$2048 \$1900 \$2104 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4916 \$16 \$2104 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4917 \$16 \$2098 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4918 \$153 \$2091 \$1900 \$2098 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4919 \$153 \$2091 \$1993 \$1771 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4920 \$16 \$2104 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4921 \$153 \$2080 \$1715 \$1674 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4923 \$153 \$2163 \$1880 \$2104 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4924 \$16 \$2098 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4925 \$153 \$2164 \$1880 \$2098 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4926 \$16 \$829 \$1929 \$2165 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$4928 \$153 \$1711 \$1928 \$2105 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4930 \$16 \$2105 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4931 \$16 \$829 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4933 \$16 \$2098 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4934 \$153 \$1992 \$1928 \$2098 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4935 \$153 \$2123 \$2092 \$1542 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4936 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$4937 \$16 \$2098 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4938 \$153 \$2051 \$1903 \$2098 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4939 \$16 \$2105 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4941 \$153 \$2052 \$1903 \$2105 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4943 \$153 \$2018 \$1854 \$2104 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4945 \$16 \$2105 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4946 \$153 \$2125 \$1854 \$2105 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4947 \$16 \$2124 \$16 \$153 \$901 VNB sky130_fd_sc_hd__clkbuf_2
X$4949 \$153 \$2125 \$2438 \$1996 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4950 \$153 \$2168 \$1782 \$1812 \$1970 \$1831 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$4951 \$153 \$1970 \$1831 \$2053 \$1782 \$1812 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$4952 \$16 \$2126 \$16 \$153 \$1782 VNB sky130_fd_sc_hd__clkbuf_2
X$4953 \$16 \$2106 \$16 \$153 \$594 VNB sky130_fd_sc_hd__clkbuf_2
X$4954 \$153 \$2106 \$1883 \$1855 \$1905 \$1971 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$4955 \$153 \$1905 \$1971 \$2107 \$1883 \$1855 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$4958 \$16 \$2107 \$16 \$153 \$964 VNB sky130_fd_sc_hd__clkbuf_2
X$4959 \$16 \$2127 \$16 \$153 \$902 VNB sky130_fd_sc_hd__clkbuf_2
X$4960 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$4962 \$16 \$964 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4963 \$153 \$2128 \$2271 \$1999 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4964 \$153 \$2082 \$1936 \$1999 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4965 \$153 \$2169 \$1906 \$2192 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4966 \$16 \$2192 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4968 \$153 \$2169 \$2269 \$1999 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4969 \$16 \$964 \$16 \$153 \$2129 VNB sky130_fd_sc_hd__inv_1
X$4970 \$16 \$964 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4972 \$153 \$2083 \$2086 \$2129 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4973 \$153 \$2170 \$1974 \$2031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4974 \$153 \$2084 \$2056 \$2129 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4975 \$16 \$2093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4976 \$16 \$354 \$1972 \$2108 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$4978 \$153 \$2057 \$1909 \$2093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4979 \$16 \$1972 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4980 \$16 \$2093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4981 \$153 \$2171 \$2058 \$2093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4982 \$16 \$354 \$16 \$153 \$2172 VNB sky130_fd_sc_hd__inv_1
X$4984 \$153 \$2094 \$2058 \$2085 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4987 \$153 \$2094 \$2271 \$2172 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4988 \$16 \$1860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4989 \$153 \$2174 \$2099 \$1973 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4990 \$153 \$2174 \$2056 \$2239 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4991 \$16 \$2093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4992 \$16 \$948 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4993 \$16 \$1885 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4994 \$16 \$608 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4995 \$16 \$1885 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$4996 \$153 \$2130 \$1936 \$2020 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$4998 \$153 \$2130 \$1886 \$2031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$4999 \$153 \$1939 \$2056 \$2020 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5000 \$153 \$2095 \$2004 \$2093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5001 \$153 \$2095 \$2265 \$1940 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5002 \$16 \$1960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5003 \$16 \$1601 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5004 \$16 \$1758 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5006 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$5007 \$16 \$2093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5008 \$153 \$2177 \$1938 \$2093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5009 \$153 \$2061 \$1938 \$2191 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5010 \$16 \$2192 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5011 \$153 \$2062 \$1938 \$2192 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5013 \$153 \$2131 \$2056 \$2032 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5015 \$153 \$2132 \$2269 \$2032 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5016 \$153 \$2133 \$1936 \$2178 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5017 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$5019 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$5020 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$5021 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$5022 \$153 \$4841 \$4864 \$3709 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5023 \$153 \$4841 \$3606 \$4859 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5024 \$16 \$3709 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5025 \$153 \$4809 \$4864 \$3473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5026 \$16 \$4902 \$16 \$153 \$4859 VNB sky130_fd_sc_hd__inv_1
X$5027 \$16 \$3473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5028 \$16 \$5152 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5030 \$16 \$4538 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5032 \$153 \$4703 \$4788 \$3615 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5033 \$16 \$3615 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5034 \$16 \$3709 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5036 \$16 \$4893 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5037 \$153 \$4704 \$4788 \$3473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5038 \$153 \$4810 \$3490 \$4692 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5039 \$16 \$3473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5040 \$16 \$3766 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5043 \$153 \$4894 \$4614 \$3385 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5044 \$16 \$3385 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5045 \$16 \$3766 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5047 \$16 \$5080 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5049 \$153 \$4895 \$4789 \$3709 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5050 \$153 \$4897 \$4789 \$3473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5052 \$16 \$3473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5053 \$16 \$3709 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5054 \$16 \$4896 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5056 \$153 \$4811 \$3307 \$4527 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5058 \$153 \$4898 \$4865 \$3766 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5059 \$16 \$3615 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5060 \$16 \$3766 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5062 \$16 \$3571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5063 \$153 \$4899 \$4865 \$3473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5065 \$153 \$4866 \$3490 \$4940 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5067 \$153 \$4900 \$4867 \$3709 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5068 \$153 \$4868 \$3478 \$4359 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5070 \$153 \$4790 \$4867 \$3474 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5071 \$16 \$3474 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5072 \$16 \$4600 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5075 \$153 \$4842 \$4791 \$3473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5076 \$153 \$4842 \$3540 \$4941 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5078 \$153 \$4843 \$4791 \$3709 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5079 \$153 \$4843 \$3606 \$4941 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5080 \$16 \$4712 \$16 \$153 \$4329 VNB sky130_fd_sc_hd__inv_1
X$5082 \$153 \$4844 \$4711 \$3709 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5083 \$153 \$4844 \$3606 \$4694 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5084 \$153 \$4746 \$3307 \$4694 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5085 \$16 \$4822 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5087 \$16 \$4860 \$16 \$153 \$4869 VNB sky130_fd_sc_hd__clkbuf_2
X$5088 \$153 \$4860 \$4715 \$4598 \$4659 \$4714 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$5089 \$16 \$4078 \$16 \$153 \$4714 VNB sky130_fd_sc_hd__clkbuf_2
X$5092 \$16 \$4747 \$16 \$153 \$4712 VNB sky130_fd_sc_hd__clkbuf_2
X$5093 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$5095 \$153 \$4793 \$4717 \$4662 \$4716 \$4661 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$5096 \$153 \$4717 \$4716 \$4901 \$4661 \$4662 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$5097 \$16 \$4662 \$4661 \$4717 \$4716 \$16 \$153 \$4870 VNB
+ sky130_fd_sc_hd__and4_2
X$5098 \$16 \$4748 \$16 \$153 \$4621 VNB sky130_fd_sc_hd__clkbuf_2
X$5099 \$16 \$4870 \$16 \$153 \$4902 VNB sky130_fd_sc_hd__clkbuf_2
X$5101 \$153 \$4815 \$3608 \$4529 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5103 \$153 \$4871 \$3608 \$4861 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5104 \$153 \$4749 \$3101 \$4529 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5105 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$5107 \$153 \$4872 \$4926 \$3620 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5108 \$153 \$4872 \$3645 \$4861 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5109 \$16 \$3620 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5110 \$16 \$3386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5113 \$153 \$4903 \$4873 \$3621 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5114 \$16 \$3621 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5115 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$5117 \$153 \$4845 \$4873 \$3620 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5118 \$153 \$4845 \$3645 \$4796 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5119 \$16 \$3620 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5120 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$5121 \$16 \$4896 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5123 \$153 \$4874 \$3435 \$4796 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5125 \$153 \$4904 \$4797 \$3620 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5126 \$153 \$4846 \$4622 \$3480 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5127 \$153 \$4846 \$3504 \$4530 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5128 \$16 \$3480 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5129 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$5131 \$16 \$3543 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5132 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$5133 \$153 \$4928 \$4875 \$3621 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5134 \$16 \$3621 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5135 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$5137 \$153 \$4862 \$4875 \$3620 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5138 \$153 \$4862 \$3645 \$4798 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5139 \$16 \$3620 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5142 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$5143 \$153 \$4905 \$4876 \$3492 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5144 \$153 \$4775 \$3504 \$4498 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5146 \$153 \$4847 \$4876 \$3620 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5147 \$153 \$4847 \$3645 \$4696 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5148 \$16 \$3620 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5151 \$153 \$4721 \$5065 \$4877 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$5152 \$16 \$3621 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5154 \$153 \$4906 \$4721 \$3621 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5155 \$153 \$4848 \$4721 \$3480 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5156 \$16 \$3480 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5157 \$16 \$3492 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5161 \$16 \$3573 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5162 \$16 \$3386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5163 \$153 \$4826 \$3354 \$4776 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5164 \$153 \$4849 \$4721 \$3386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5165 \$153 \$4849 \$3435 \$4776 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5166 \$153 \$4907 \$4799 \$3960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5168 \$153 \$4863 \$3079 \$5066 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5169 \$16 \$3960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5170 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$5171 \$16 \$3791 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5172 \$153 \$4850 \$4799 \$3791 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5173 \$153 \$4850 \$3919 \$4801 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5175 \$16 \$3792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5176 \$16 \$3791 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5178 \$153 \$4754 \$3716 \$4697 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5180 \$153 \$4722 \$4759 \$4878 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$5181 \$153 \$4851 \$4722 \$4048 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5182 \$153 \$4851 \$3858 \$4697 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5184 \$153 \$4852 \$4698 \$3960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5186 \$153 \$4879 \$3919 \$4637 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5187 \$153 \$4880 \$4698 \$3889 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5188 \$16 \$4475 \$16 \$153 \$4881 VNB sky130_fd_sc_hd__clkbuf_2
X$5189 \$16 \$3889 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5190 \$16 \$3852 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5191 \$153 \$4853 \$4638 \$3852 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5192 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$5194 \$16 \$3960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5196 \$153 \$4854 \$4638 \$3960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5197 \$153 \$4908 \$4638 \$3792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5198 \$16 \$4562 \$4724 \$4725 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$5199 \$16 \$4882 \$16 \$153 \$4587 VNB sky130_fd_sc_hd__inv_1
X$5200 \$153 \$4909 \$4726 \$3889 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5202 \$153 \$4910 \$4726 \$3792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5203 \$16 \$4837 \$4724 \$4828 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$5205 \$153 \$4883 \$4726 \$3960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5206 \$153 \$4728 \$3763 \$4639 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5207 \$153 \$4883 \$3716 \$4639 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5209 \$153 \$4911 \$4804 \$3960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5210 \$16 \$3960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5212 \$153 \$4729 \$4804 \$3731 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5213 \$16 \$4048 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5214 \$153 \$4884 \$4804 \$3814 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5215 \$16 \$4830 \$16 \$153 \$4700 VNB sky130_fd_sc_hd__inv_1
X$5217 \$153 \$4832 \$3919 \$4700 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5218 \$153 \$4884 \$3651 \$4700 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5219 \$16 \$4305 \$16 \$153 \$4912 VNB sky130_fd_sc_hd__clkbuf_2
X$5220 \$16 \$4834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5221 \$153 \$4461 \$3676 \$5158 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5222 \$153 \$4782 \$4414 \$4954 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5223 \$153 \$4731 \$4759 \$4886 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$5225 \$153 \$4806 \$4887 \$3898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5226 \$16 \$4930 \$16 \$153 \$4643 VNB sky130_fd_sc_hd__inv_1
X$5227 \$153 \$4888 \$4887 \$4057 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5228 \$16 \$4569 \$16 \$153 \$4958 VNB sky130_fd_sc_hd__clkbuf_2
X$5230 \$153 \$4855 \$4887 \$3680 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5232 \$16 \$4129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5234 \$153 \$4855 \$3719 \$4807 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5235 \$16 \$3680 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5236 \$16 \$3602 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5238 \$153 \$4913 \$4626 \$3898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5240 \$16 \$4129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5241 \$16 \$4613 \$16 \$153 \$5116 VNB sky130_fd_sc_hd__clkbuf_2
X$5242 \$153 \$4856 \$4626 \$4129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5245 \$153 \$4856 \$3986 \$4484 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5247 \$153 \$4206 \$3986 \$4379 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5248 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$5249 \$153 \$4889 \$3676 \$4808 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5250 \$153 \$5076 \$3719 \$4808 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5251 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$5252 \$16 \$4882 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5253 \$153 \$4890 \$3860 \$4808 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5255 \$153 \$4923 \$3565 \$4808 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5256 \$153 \$4284 \$3860 \$4379 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5257 \$153 \$4285 \$4414 \$4379 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5259 \$16 \$4837 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5260 \$153 \$4591 \$3986 \$4857 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5261 \$153 \$4286 \$3676 \$4857 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5262 \$16 \$4837 \$4736 \$4914 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$5263 \$16 \$4129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5266 \$153 \$4915 \$4739 \$3721 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5267 \$16 \$4837 \$16 \$153 \$4646 VNB sky130_fd_sc_hd__inv_1
X$5268 \$16 \$3721 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5269 \$153 \$4858 \$4739 \$3602 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5270 \$153 \$4891 \$3719 \$4646 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5271 \$153 \$4858 \$3565 \$4646 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5274 \$16 \$3602 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5275 \$153 \$5098 \$4892 \$3602 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5276 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$5277 \$153 \$4593 \$3565 \$4537 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5278 \$153 \$4916 \$4740 \$3898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5279 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$5282 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$5283 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$5284 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$5285 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$5286 \$153 \$4925 \$4864 \$3474 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5287 \$16 \$3474 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5288 \$16 \$3766 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5289 \$16 \$4902 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5291 \$153 \$4925 \$3490 \$4859 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5293 \$153 \$4968 \$4864 \$3615 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5294 \$16 \$3615 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5295 \$153 \$4917 \$4788 \$3616 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5296 \$153 \$4917 \$3389 \$4692 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5297 \$16 \$3616 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5300 \$16 \$4893 \$16 \$153 \$4692 VNB sky130_fd_sc_hd__inv_1
X$5301 \$153 \$4969 \$4788 \$3766 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5302 \$16 \$3385 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5304 \$153 \$4970 \$4614 \$3766 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5305 \$153 \$4970 \$3478 \$4707 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5306 \$153 \$5535 \$5107 \$4579 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5308 \$153 \$4708 \$4789 \$3474 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5309 \$16 \$3474 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5310 \$153 \$4971 \$4789 \$3766 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5311 \$16 \$3766 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5313 \$16 \$4939 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5314 \$153 \$4972 \$4865 \$3709 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5317 \$16 \$3709 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5319 \$153 \$4898 \$3478 \$4940 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5320 \$153 \$4866 \$4865 \$3474 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5321 \$16 \$3474 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5322 \$16 \$3473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5323 \$16 \$4973 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5325 \$153 \$4868 \$4867 \$3766 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5326 \$16 \$3766 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5328 \$16 \$3709 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5330 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$5331 \$153 \$4786 \$4867 \$3473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5332 \$16 \$3473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5334 \$16 \$5026 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5335 \$16 \$3615 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5336 \$153 \$4974 \$4791 \$3615 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5337 \$153 \$4974 \$3307 \$4941 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5338 \$16 \$3473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5340 \$153 \$4814 \$3490 \$4941 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5341 \$16 \$3385 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5343 \$16 \$4869 \$4012 \$4975 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$5344 \$16 \$3571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5345 \$16 \$3385 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5346 \$153 \$4942 \$4711 \$3385 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5347 \$153 \$4942 \$3394 \$4694 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5349 \$16 \$4822 \$16 \$153 \$4694 VNB sky130_fd_sc_hd__inv_1
X$5350 \$16 \$3709 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5351 \$16 \$4712 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5352 \$16 \$4943 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5354 \$153 \$4944 \$3478 \$4694 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5355 \$16 \$4945 \$16 \$153 \$3907 VNB sky130_fd_sc_hd__clkbuf_2
X$5356 \$153 \$4976 \$4659 \$4598 \$4715 \$4714 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$5357 \$153 \$4945 \$4714 \$4598 \$4659 \$4715 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$5358 \$16 \$4946 \$16 \$153 \$4494 VNB sky130_fd_sc_hd__clkbuf_2
X$5360 \$16 \$4079 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5361 \$153 \$4977 \$4716 \$4717 \$4661 \$4662 \$16 \$16 VNB
+ sky130_fd_sc_hd__nor4b_2
X$5362 \$16 \$4901 \$16 \$153 \$5080 VNB sky130_fd_sc_hd__clkbuf_2
X$5364 \$153 \$4717 \$4661 \$4978 \$4716 \$4662 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$5366 \$153 \$4871 \$4926 \$3621 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5368 \$153 \$4918 \$4926 \$3573 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5369 \$153 \$4918 \$3079 \$4861 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5370 \$16 \$3573 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5373 \$153 \$4980 \$4926 \$3386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5374 \$153 \$4980 \$3435 \$4861 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5376 \$153 \$4795 \$4873 \$3573 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5377 \$153 \$4903 \$3608 \$4796 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5378 \$16 \$3573 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5379 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$5381 \$153 \$4874 \$4873 \$3386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5382 \$16 \$3386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5383 \$153 \$4817 \$4797 \$3386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5384 \$16 \$3386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5386 \$16 \$3573 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5388 \$153 \$4819 \$4797 \$3621 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5390 \$153 \$4904 \$3645 \$4818 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5391 \$153 \$4927 \$3556 \$4818 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5392 \$16 \$4947 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5393 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$5394 \$153 \$4820 \$4875 \$3573 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5395 \$16 \$3573 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5396 \$153 \$4928 \$3608 \$4798 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5399 \$153 \$4919 \$4875 \$3386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5400 \$153 \$4919 \$3435 \$4798 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5401 \$16 \$3386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5403 \$16 \$3573 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5404 \$153 \$4981 \$4876 \$3573 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5405 \$153 \$4669 \$3354 \$4498 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5407 \$153 \$4823 \$4876 \$3621 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5408 \$16 \$3621 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5410 \$16 \$4712 \$3957 \$4877 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$5411 \$153 \$4982 \$4948 \$3621 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5412 \$153 \$4825 \$4948 \$3620 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5414 \$16 \$3620 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5415 \$16 \$3480 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5416 \$153 \$4906 \$3608 \$4776 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5417 \$16 \$3621 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5418 \$16 \$4712 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5420 \$153 \$4984 \$4948 \$3386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5421 \$153 \$4863 \$4948 \$3573 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5422 \$16 \$3386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5423 \$16 \$5209 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5424 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5426 \$153 \$3822 \$1482 \$5209 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5427 \$153 \$4800 \$4799 \$3889 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5428 \$153 \$4907 \$3716 \$4801 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5429 \$153 \$4929 \$3939 \$4801 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5430 \$16 \$3792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5431 \$16 \$4760 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5432 \$16 \$3852 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5434 \$153 \$4985 \$4799 \$3852 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5435 \$153 \$4986 \$4722 \$3792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5437 \$16 \$4930 \$4881 \$4878 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$5438 \$16 \$3889 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5439 \$153 \$4987 \$4722 \$3889 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5441 \$153 \$4987 \$3962 \$4697 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5442 \$16 \$4930 \$16 \$153 \$4697 VNB sky130_fd_sc_hd__inv_1
X$5444 \$153 \$4879 \$4698 \$3791 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5445 \$153 \$4698 \$4756 \$4989 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$5447 \$16 \$4949 \$16 \$153 \$4637 VNB sky130_fd_sc_hd__inv_1
X$5448 \$153 \$4950 \$3939 \$4637 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5450 \$153 \$4880 \$3962 \$4637 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5451 \$153 \$5088 \$3788 \$4951 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5453 \$153 \$4991 \$4931 \$3731 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5455 \$16 \$4562 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5456 \$16 \$3731 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5457 \$16 \$3792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5458 \$153 \$4638 \$4781 \$4932 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$5460 \$153 \$4993 \$4952 \$3731 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5461 \$16 \$3889 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5463 \$153 \$4909 \$3962 \$4639 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5464 \$153 \$4994 \$4920 \$3731 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5465 \$153 \$4994 \$3788 \$4953 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5466 \$16 \$4837 \$16 \$153 \$4639 VNB sky130_fd_sc_hd__inv_1
X$5468 \$153 \$4996 \$5043 \$3731 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5470 \$16 \$4997 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5471 \$16 \$4954 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5472 \$16 \$3889 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5473 \$153 \$4999 \$4804 \$3889 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5474 \$16 \$4724 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5475 \$153 \$5073 \$3763 \$4700 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5476 \$16 \$4830 \$4724 \$5000 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$5479 \$153 \$4911 \$3716 \$4700 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5480 \$153 \$4783 \$3939 \$4700 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5482 \$153 \$4955 \$3858 \$4700 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5483 \$16 \$4956 \$16 \$153 \$4930 VNB sky130_fd_sc_hd__clkbuf_2
X$5484 \$16 \$4317 \$16 \$153 \$4933 VNB sky130_fd_sc_hd__clkbuf_2
X$5485 \$153 \$4934 \$4933 \$4912 \$4833 \$4935 \$16 \$16 VNB
+ sky130_fd_sc_hd__nor4b_2
X$5486 \$16 \$4958 \$4937 \$4936 \$5001 \$16 \$153 \$4957 VNB
+ sky130_fd_sc_hd__and4_2
X$5488 \$16 \$4934 \$16 \$153 \$4949 VNB sky130_fd_sc_hd__clkbuf_2
X$5490 \$153 \$4921 \$5001 \$4958 \$4936 \$4937 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$5491 \$153 \$4938 \$4937 \$4958 \$4936 \$5001 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$5492 \$153 \$4959 \$4887 \$3826 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5493 \$153 \$4959 \$3893 \$4807 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5494 \$16 \$4305 \$16 \$153 \$4936 VNB sky130_fd_sc_hd__clkbuf_2
X$5495 \$16 \$3721 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5497 \$16 \$3898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5499 \$153 \$5004 \$3142 \$4807 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5500 \$153 \$4922 \$4887 \$4129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5501 \$153 \$4960 \$4887 \$3602 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5502 \$153 \$4961 \$4414 \$5019 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5504 \$16 \$4949 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5507 \$16 \$3826 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5508 \$153 \$4962 \$3142 \$4484 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5510 \$153 \$5005 \$4626 \$3826 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5511 \$16 \$4963 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5512 \$16 \$4963 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5513 \$16 \$4964 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5514 \$16 \$3721 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5515 \$153 \$4889 \$4627 \$3721 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5516 \$16 \$4949 \$16 \$153 \$4808 VNB sky130_fd_sc_hd__inv_1
X$5519 \$16 \$3602 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5520 \$153 \$4923 \$4627 \$3602 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5521 \$16 \$4781 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5522 \$153 \$4737 \$4781 \$5006 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$5523 \$153 \$4924 \$4737 \$3680 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5524 \$16 \$4882 \$16 \$153 \$3567 VNB sky130_fd_sc_hd__inv_1
X$5525 \$16 \$3826 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5527 \$153 \$5007 \$4737 \$3826 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5528 \$153 \$4739 \$4803 \$4914 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$5529 \$153 \$5008 \$4739 \$3691 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5530 \$153 \$4763 \$3893 \$4646 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5533 \$153 \$4891 \$4739 \$3680 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5534 \$16 \$4830 \$4736 \$5009 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$5536 \$16 \$4129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5537 \$153 \$5010 \$4892 \$4129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5538 \$16 \$4830 \$16 \$153 \$5011 VNB sky130_fd_sc_hd__inv_1
X$5539 \$16 \$4830 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5541 \$153 \$4966 \$3565 \$4965 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5543 \$16 \$4057 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5544 \$16 \$3898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5545 \$153 \$5510 \$4740 \$4057 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5547 \$153 \$4594 \$3676 \$4537 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5548 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$5549 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$5550 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$5551 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$5553 \$153 \$4242 \$4241 \$3709 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5554 \$153 \$4382 \$3389 \$4372 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5555 \$16 \$3709 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5557 \$153 \$4416 \$4241 \$3473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5558 \$16 \$3473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5559 \$16 \$5376 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5562 \$153 \$4470 \$4241 \$3615 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5563 \$16 \$4320 \$16 \$153 \$4066 VNB sky130_fd_sc_hd__inv_1
X$5565 \$153 \$4417 \$4158 \$3474 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5566 \$16 \$3474 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5567 \$16 \$3766 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5568 \$153 \$4418 \$4383 \$3616 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5570 \$16 \$3616 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5572 \$153 \$4326 \$3540 \$4067 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5573 \$16 \$3473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5575 \$153 \$4327 \$3394 \$4067 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5576 \$16 \$3571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5577 \$16 \$3385 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5578 \$16 \$4178 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5579 \$153 \$4384 \$3422 \$4489 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5581 \$153 \$4358 \$4143 \$3616 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5583 \$16 \$3616 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5584 \$16 \$3615 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5586 \$153 \$4358 \$3389 \$4328 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5588 \$153 \$4419 \$4143 \$3474 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5589 \$153 \$4143 \$5388 \$4385 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$5590 \$16 \$4181 \$16 \$153 \$4538 VNB sky130_fd_sc_hd__clkbuf_2
X$5591 \$16 \$4421 \$16 \$153 \$4328 VNB sky130_fd_sc_hd__inv_1
X$5592 \$16 \$3571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5593 \$16 \$5388 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5595 \$153 \$4420 \$4386 \$3616 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5596 \$153 \$4387 \$3540 \$4373 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5598 \$153 \$4388 \$3307 \$4359 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5600 \$153 \$4389 \$3606 \$4373 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5601 \$16 \$4181 \$16 \$153 \$4012 VNB sky130_fd_sc_hd__clkbuf_2
X$5602 \$16 \$5125 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5603 \$16 \$5349 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5605 \$16 \$2743 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5607 \$153 \$4391 \$4390 \$3766 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5608 \$153 \$4391 \$3478 \$4329 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5609 \$153 \$4245 \$4319 \$3385 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5610 \$153 \$4446 \$3478 \$4230 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5611 \$16 \$3385 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5612 \$16 \$3766 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5613 \$16 \$3473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5615 \$153 \$4422 \$4319 \$3473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5616 \$153 \$4133 \$3389 \$4019 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5617 \$153 \$4331 \$3606 \$4230 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5618 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$5619 \$16 \$4620 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5620 \$16 \$4472 \$16 \$153 \$4106 VNB sky130_fd_sc_hd__clkbuf_2
X$5621 \$153 \$4374 \$4393 \$4394 \$4392 \$4447 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$5623 \$16 \$4360 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5626 \$16 \$4360 \$16 \$153 \$2387 VNB sky130_fd_sc_hd__clkbuf_2
X$5627 \$16 \$4395 \$16 \$153 \$4421 VNB sky130_fd_sc_hd__clkbuf_2
X$5628 \$16 \$4394 \$16 \$153 \$3997 VNB sky130_fd_sc_hd__clkbuf_2
X$5629 \$16 \$3911 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5630 \$16 \$4215 \$4110 \$4148 \$4160 \$16 \$153 \$4423 VNB
+ sky130_fd_sc_hd__and4_2
X$5632 \$16 \$4275 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5633 \$16 \$4320 \$4275 \$4396 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$5634 \$16 \$4397 \$16 \$153 \$4215 VNB sky130_fd_sc_hd__clkbuf_2
X$5636 \$153 \$4424 \$4321 \$3572 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5637 \$16 \$4320 \$16 \$153 \$4216 VNB sky130_fd_sc_hd__inv_1
X$5640 \$16 \$3572 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5642 \$153 \$4425 \$4321 \$3543 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5643 \$153 \$4361 \$4321 \$3480 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5644 \$153 \$4336 \$4321 \$3386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5645 \$16 \$3480 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5646 \$16 \$3386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5650 \$153 \$3954 \$4179 \$4273 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$5651 \$16 \$4178 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5652 \$153 \$4522 \$3354 \$4633 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5653 \$16 \$3572 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5654 \$16 \$4269 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5656 \$153 \$4362 \$4398 \$3620 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5657 \$153 \$4362 \$3645 \$4338 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5659 \$153 \$4473 \$4398 \$3621 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5660 \$153 \$4322 \$5388 \$4399 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$5662 \$153 \$4250 \$4322 \$3573 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5663 \$153 \$4523 \$3556 \$4300 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5666 \$153 \$4251 \$4322 \$3492 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5667 \$16 \$3492 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5669 \$16 \$4106 \$4014 \$4400 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$5670 \$153 \$4163 \$5125 \$4400 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$5672 \$153 \$4426 \$4163 \$3572 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5674 \$16 \$4106 \$16 \$153 \$4164 VNB sky130_fd_sc_hd__inv_1
X$5675 \$16 \$3572 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5676 \$16 \$3543 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5678 \$153 \$4375 \$4163 \$3492 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5679 \$153 \$4375 \$3354 \$4164 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5680 \$153 \$4427 \$3079 \$4164 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5681 \$16 \$4246 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5682 \$16 \$4340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5683 \$153 \$4401 \$3504 \$4363 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5686 \$153 \$4402 \$3435 \$4363 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5687 \$153 \$4403 \$3354 \$4363 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5689 \$153 \$4342 \$4194 \$3621 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5690 \$16 \$3621 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5692 \$153 \$4428 \$4404 \$3480 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5693 \$16 \$3480 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5695 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$5696 \$153 \$153 \$3354 \$4233 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5697 \$16 \$3386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5698 \$153 \$4364 \$4404 \$3386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5699 \$153 \$4364 \$3435 \$4501 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5700 \$16 \$3543 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5702 \$16 \$3272 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5703 \$16 \$3916 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5704 \$16 \$3983 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5705 \$16 \$3763 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5706 \$16 \$3814 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5707 \$16 \$3889 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5708 \$16 \$3960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5710 \$153 \$4429 \$4481 \$3814 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5712 \$153 \$4365 \$4254 \$4048 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5713 \$153 \$4365 \$3858 \$4234 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5714 \$153 \$4343 \$3962 \$4234 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5715 \$16 \$4324 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5717 \$16 \$4324 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5719 \$16 \$3731 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5721 \$16 \$4324 \$16 \$153 \$4234 VNB sky130_fd_sc_hd__inv_1
X$5722 \$16 \$4430 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5723 \$153 \$4405 \$3716 \$4234 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5724 \$153 \$4431 \$3788 \$4234 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5725 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$5727 \$153 \$4278 \$3919 \$4235 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5728 \$153 \$4406 \$3962 \$4235 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5729 \$16 \$4432 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5730 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$5731 \$16 \$3814 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5734 \$16 \$3792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5735 \$153 \$4407 \$3939 \$4235 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5736 \$16 \$3960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5738 \$153 \$4151 \$4256 \$3814 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5739 \$16 \$3889 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5740 \$16 \$4415 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5742 \$16 \$4048 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5743 \$153 \$4474 \$4256 \$4048 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5744 \$16 \$3792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5746 \$16 \$4415 \$16 \$153 \$4167 VNB sky130_fd_sc_hd__inv_1
X$5747 \$153 \$4433 \$4257 \$3792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5748 \$153 \$4302 \$3788 \$4167 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5750 \$16 \$3852 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5751 \$153 \$4476 \$4257 \$3852 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5752 \$153 \$4346 \$3858 \$4509 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5754 \$153 \$4366 \$4323 \$3791 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5755 \$153 \$4366 \$3919 \$4236 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5756 \$153 \$4434 \$4323 \$3731 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5757 \$153 \$4409 \$3858 \$4236 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5758 \$16 \$4464 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5759 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$5761 \$16 \$3852 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5762 \$153 \$4201 \$3962 \$4024 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5763 \$153 \$4435 \$4260 \$3852 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5765 \$16 \$4048 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5766 \$153 \$4367 \$4260 \$4048 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5767 \$153 \$4367 \$3858 \$4237 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5770 \$153 \$4260 \$4316 \$4463 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$5771 \$16 \$2936 \$16 \$153 \$4347 VNB sky130_fd_sc_hd__clkbuf_2
X$5772 \$16 \$2793 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5773 \$16 \$3983 \$16 \$153 \$4436 VNB sky130_fd_sc_hd__clkbuf_2
X$5774 \$16 \$4376 \$16 \$153 \$4237 VNB sky130_fd_sc_hd__inv_1
X$5775 \$16 \$4317 \$16 \$153 \$4265 VNB sky130_fd_sc_hd__clkbuf_2
X$5776 \$16 \$4305 \$16 \$153 \$4239 VNB sky130_fd_sc_hd__clkbuf_2
X$5777 \$16 \$2936 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5778 \$153 \$4377 \$4265 \$4239 \$4266 \$4225 \$16 \$16 VNB
+ sky130_fd_sc_hd__nor4b_2
X$5779 \$16 \$4377 \$16 \$153 \$4376 VNB sky130_fd_sc_hd__clkbuf_2
X$5781 \$16 \$3898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5783 \$16 \$4324 \$3988 \$4437 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$5784 \$16 \$4780 \$3988 \$4438 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$5785 \$16 \$4349 \$16 \$153 \$4464 VNB sky130_fd_sc_hd__clkbuf_2
X$5787 \$153 \$4410 \$3860 \$3567 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5788 \$153 \$3827 \$3565 \$3461 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5789 \$153 \$4411 \$4414 \$4378 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5790 \$16 \$4780 \$16 \$153 \$4378 VNB sky130_fd_sc_hd__inv_1
X$5791 \$16 \$3680 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5792 \$153 \$4368 \$3142 \$4378 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5794 \$153 \$4368 \$4483 \$3691 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5795 \$16 \$3691 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5797 \$16 \$3602 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5798 \$153 \$4413 \$4483 \$3602 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5799 \$153 \$4412 \$3986 \$4378 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5800 \$153 \$4413 \$3565 \$4378 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5803 \$153 \$4059 \$4414 \$3895 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5804 \$16 \$4415 \$3988 \$4439 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$5805 \$16 \$4415 \$16 \$153 \$4379 VNB sky130_fd_sc_hd__inv_1
X$5806 \$153 \$4440 \$4095 \$3691 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5807 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$5808 \$16 \$3826 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5809 \$153 \$4370 \$4325 \$3826 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5812 \$153 \$4370 \$3893 \$4369 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5813 \$153 \$4351 \$3565 \$4369 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5814 \$153 \$4207 \$3676 \$4379 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5815 \$153 \$4440 \$3142 \$4379 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5816 \$153 \$4318 \$3719 \$4379 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5817 \$16 \$4562 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5818 \$153 \$4288 \$3676 \$4371 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5820 \$16 \$3898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5822 \$16 \$4464 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5823 \$16 \$4464 \$16 \$153 \$4371 VNB sky130_fd_sc_hd__inv_1
X$5824 \$153 \$4380 \$4414 \$4171 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5825 \$153 \$3614 \$3565 \$4171 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5826 \$153 \$3759 \$3142 \$4171 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5827 \$153 \$4172 \$4316 \$4381 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$5828 \$16 \$4376 \$4156 \$4381 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$5829 \$16 \$3691 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5831 \$153 \$4356 \$4172 \$3680 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5832 \$16 \$4376 \$16 \$153 \$4173 VNB sky130_fd_sc_hd__inv_1
X$5833 \$16 \$4376 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5834 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$5835 \$153 \$4291 \$3565 \$4173 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5836 \$16 \$4057 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5837 \$153 \$4098 \$4172 \$4057 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5838 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$5841 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$5842 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$5843 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$5844 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$5846 \$153 \$4441 \$4241 \$3474 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5847 \$16 \$3474 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5848 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$5851 \$153 \$4241 \$5376 \$4486 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$5852 \$153 \$4487 \$4469 \$3615 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5853 \$153 \$4416 \$3540 \$4066 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5854 \$153 \$4470 \$3307 \$4066 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5855 \$16 \$3615 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5856 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$5859 \$16 \$3474 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5860 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$5861 \$153 \$4488 \$4383 \$3766 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5862 \$16 \$3473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5863 \$16 \$3766 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5865 \$153 \$4442 \$4383 \$3385 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5866 \$153 \$4442 \$3394 \$4489 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5867 \$16 \$3385 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5869 \$153 \$4471 \$3606 \$4489 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5870 \$16 \$4479 \$16 \$153 \$4489 VNB sky130_fd_sc_hd__inv_1
X$5871 \$16 \$3709 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5872 \$153 \$4443 \$4143 \$3615 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5873 \$153 \$4444 \$4617 \$3474 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5874 \$153 \$4443 \$3307 \$4328 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5878 \$16 \$3474 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5879 \$153 \$4419 \$3490 \$4328 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5880 \$16 \$4421 \$4144 \$4385 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$5881 \$16 \$4621 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5882 \$16 \$4421 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5884 \$16 \$4421 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5885 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$5887 \$153 \$4445 \$4386 \$3474 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5888 \$153 \$4445 \$3490 \$4373 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5891 \$153 \$4490 \$4386 \$3766 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5892 \$16 \$3766 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5894 \$153 \$4491 \$4390 \$3709 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5895 \$153 \$4330 \$4390 \$3616 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5896 \$16 \$3616 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5897 \$16 \$3709 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5899 \$153 \$4446 \$4319 \$3766 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5900 \$153 \$4492 \$3307 \$4329 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5901 \$153 \$4493 \$3307 \$4230 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5902 \$153 \$4332 \$4319 \$3616 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5903 \$16 \$3616 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5904 \$16 \$4494 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5907 \$16 \$4495 \$16 \$153 \$4178 VNB sky130_fd_sc_hd__clkbuf_2
X$5908 \$16 \$4619 \$16 \$153 \$4229 VNB sky130_fd_sc_hd__clkbuf_2
X$5909 \$153 \$4472 \$4392 \$4374 \$4393 \$4447 \$16 \$16 VNB
+ sky130_fd_sc_hd__nor4b_2
X$5910 \$153 \$4392 \$4393 \$4395 \$4374 \$4447 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$5911 \$16 \$4272 \$16 \$153 \$4374 VNB sky130_fd_sc_hd__clkbuf_2
X$5913 \$16 \$2387 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5914 \$16 \$2387 \$16 \$153 \$4496 VNB sky130_fd_sc_hd__clkbuf_2
X$5915 \$16 \$4496 \$4539 \$4497 \$153 \$4397 \$16 VNB sky130_fd_sc_hd__and3b_4
X$5916 \$16 \$2233 \$16 \$153 \$4497 VNB sky130_fd_sc_hd__clkbuf_2
X$5917 \$16 \$2233 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5919 \$153 \$4321 \$5376 \$4396 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$5920 \$16 \$5376 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5921 \$16 \$4039 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5923 \$16 \$4320 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5924 \$153 \$4335 \$3608 \$4216 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5925 \$153 \$4424 \$3101 \$4216 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5926 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$5927 \$153 \$4425 \$3556 \$4216 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5928 \$16 \$3543 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5931 \$153 \$4448 \$4321 \$3620 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5932 \$153 \$4448 \$3645 \$4216 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5933 \$16 \$3620 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5935 \$153 \$4449 \$4540 \$3480 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5936 \$153 \$4449 \$3504 \$4633 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5940 \$153 \$4337 \$4398 \$3573 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5942 \$16 \$3620 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5943 \$16 \$3573 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5944 \$153 \$4450 \$4398 \$3386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5946 \$153 \$4473 \$3608 \$4338 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5947 \$16 \$4421 \$4014 \$4399 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$5949 \$16 \$3572 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5952 \$153 \$4451 \$4322 \$3572 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5953 \$153 \$4451 \$3101 \$4300 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5955 \$153 \$4452 \$4322 \$3620 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5956 \$153 \$4452 \$3645 \$4300 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5957 \$16 \$3620 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5958 \$16 \$5125 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5960 \$16 \$3573 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5961 \$153 \$4499 \$3079 \$4498 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5962 \$153 \$4453 \$4163 \$3543 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5963 \$153 \$4426 \$3101 \$4164 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5965 \$153 \$4427 \$4163 \$3573 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5966 \$16 \$3492 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5969 \$16 \$3573 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5971 \$153 \$4401 \$4480 \$3480 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5973 \$153 \$4500 \$3645 \$4363 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5974 \$16 \$3480 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5975 \$153 \$4454 \$4480 \$3621 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5976 \$153 \$4454 \$3608 \$4363 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5979 \$153 \$4455 \$4404 \$3572 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5980 \$153 \$4455 \$3101 \$4501 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5981 \$153 \$4428 \$3504 \$4501 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5982 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$5983 \$16 \$3620 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5984 \$153 \$4456 \$4404 \$3543 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5987 \$153 \$4456 \$3556 \$4501 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5988 \$16 \$3310 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5990 \$153 \$4502 \$4481 \$3960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5991 \$153 \$4457 \$4481 \$3889 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5992 \$16 \$4048 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5993 \$153 \$4503 \$3763 \$4531 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$5995 \$153 \$4504 \$4254 \$3792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$5996 \$16 \$4324 \$4166 \$4505 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$5997 \$16 \$3960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$5998 \$153 \$4405 \$4254 \$3960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6000 \$153 \$4406 \$4165 \$3889 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6002 \$16 \$3889 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6003 \$153 \$4506 \$3858 \$4235 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6004 \$16 \$3960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6005 \$16 \$4432 \$4166 \$4507 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$6006 \$153 \$4508 \$4165 \$3960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6007 \$153 \$4407 \$4165 \$3792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6008 \$16 \$4415 \$4166 \$4525 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$6011 \$153 \$4344 \$4256 \$3889 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6012 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$6013 \$16 \$3960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6014 \$153 \$4474 \$3858 \$4167 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6015 \$153 \$4458 \$4257 \$3960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6016 \$153 \$4458 \$3716 \$4509 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6018 \$153 \$4433 \$3939 \$4509 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6019 \$16 \$4475 \$16 \$153 \$4015 VNB sky130_fd_sc_hd__clkbuf_2
X$6021 \$153 \$4476 \$3763 \$4509 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6023 \$16 \$3791 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6024 \$153 \$4459 \$4323 \$3960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6025 \$153 \$4459 \$3716 \$4236 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6026 \$16 \$4464 \$4015 \$4510 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$6028 \$153 \$4409 \$4323 \$4048 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6029 \$16 \$4464 \$16 \$153 \$4236 VNB sky130_fd_sc_hd__inv_1
X$6030 \$16 \$5381 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6032 \$16 \$3792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6033 \$153 \$4460 \$4260 \$3792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6034 \$153 \$4460 \$3939 \$4237 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6036 \$16 \$4461 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6037 \$16 \$4376 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6038 \$16 \$3791 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6040 \$153 \$4435 \$3763 \$4237 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6041 \$153 \$4462 \$4260 \$3791 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6042 \$153 \$4462 \$3919 \$4237 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6043 \$16 \$4376 \$4015 \$4463 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$6044 \$16 \$2576 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6045 \$16 \$2233 \$16 \$153 \$4477 VNB sky130_fd_sc_hd__clkbuf_2
X$6047 \$16 \$4544 \$4436 \$4477 \$153 \$4511 \$16 VNB sky130_fd_sc_hd__and3b_4
X$6049 \$16 \$4477 \$4436 \$4544 \$153 \$4482 \$16 VNB sky130_fd_sc_hd__and3b_4
X$6050 \$153 \$4265 \$4266 \$4512 \$4239 \$4225 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$6051 \$16 \$4482 \$16 \$153 \$4225 VNB sky130_fd_sc_hd__clkbuf_2
X$6052 \$16 \$4376 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6054 \$153 \$4094 \$4430 \$4437 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$6055 \$153 \$4411 \$4483 \$4057 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6057 \$153 \$4478 \$4483 \$3826 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6058 \$153 \$4478 \$3893 \$4378 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6060 \$153 \$4465 \$4483 \$3898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6061 \$153 \$4513 \$3565 \$4643 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6062 \$16 \$4590 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6064 \$16 \$4129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6066 \$153 \$4412 \$4483 \$4129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6067 \$153 \$4095 \$4542 \$4439 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$6068 \$16 \$4432 \$3988 \$4514 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$6069 \$16 \$3691 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6070 \$153 \$4515 \$4325 \$3691 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6071 \$16 \$4432 \$16 \$153 \$4369 VNB sky130_fd_sc_hd__inv_1
X$6073 \$16 \$4432 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6074 \$16 \$4432 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6076 \$16 \$4129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6077 \$153 \$4466 \$4325 \$4129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6079 \$153 \$4466 \$3986 \$4369 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6081 \$16 \$3602 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6082 \$16 \$4129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6083 \$153 \$4516 \$4267 \$3602 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6085 \$153 \$4517 \$4267 \$3826 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6086 \$16 \$3826 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6087 \$16 \$4464 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6088 \$153 \$4467 \$3860 \$4371 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6089 \$153 \$4467 \$4268 \$3898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6090 \$16 \$3826 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6091 \$153 \$3684 \$3860 \$4171 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6093 \$153 \$4518 \$4268 \$3826 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6095 \$153 \$4519 \$4485 \$4129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6096 \$153 \$4468 \$4485 \$3691 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6097 \$16 \$4567 \$16 \$153 \$4537 VNB sky130_fd_sc_hd__inv_1
X$6098 \$16 \$4567 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6099 \$16 \$3826 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6101 \$153 \$4520 \$4485 \$3826 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6102 \$153 \$4521 \$4485 \$3898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6104 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$6105 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$6106 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$6107 \$153 \$4075 \$4241 \$3616 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6108 \$16 \$3616 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6109 \$153 \$4242 \$3606 \$4066 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6110 \$153 \$4210 \$4241 \$3385 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6111 \$16 \$3385 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6112 \$16 \$3385 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6113 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$6115 \$153 \$4175 \$3394 \$3765 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6116 \$153 \$4100 \$3307 \$3765 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6117 \$16 \$4083 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6119 \$153 \$4076 \$4158 \$3616 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6120 \$153 \$4243 \$3478 \$4067 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6121 \$153 \$4176 \$3606 \$4067 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6124 \$153 \$4177 \$4158 \$3571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6125 \$16 \$3616 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6126 \$16 \$4178 \$4144 \$4228 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$6127 \$153 \$3864 \$4269 \$4228 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$6128 \$16 \$4269 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6130 \$153 \$4270 \$4143 \$3385 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6132 \$16 \$3385 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6133 \$16 \$4229 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6135 \$153 \$4180 \$3540 \$4328 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6136 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$6137 \$153 \$4211 \$4143 \$3766 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6138 \$153 \$4211 \$3478 \$4328 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6139 \$153 \$4030 \$3307 \$3872 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6141 \$153 \$4244 \$3394 \$3875 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6142 \$153 \$4212 \$3947 \$3766 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6143 \$153 \$4212 \$3478 \$3875 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6144 \$16 \$4146 \$4144 \$4271 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$6146 \$153 \$4213 \$3838 \$3616 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6148 \$153 \$4182 \$3838 \$3766 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6149 \$16 \$4146 \$16 \$153 \$3935 VNB sky130_fd_sc_hd__inv_1
X$6150 \$16 \$3766 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6151 \$153 \$4214 \$4077 \$3571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6152 \$153 \$4214 \$3422 \$4019 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6153 \$153 \$4245 \$3394 \$4230 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6156 \$16 \$3474 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6157 \$16 \$2634 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6158 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$6159 \$153 \$4077 \$4246 \$4109 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$6160 \$16 \$3886 \$16 \$153 \$4019 VNB sky130_fd_sc_hd__inv_1
X$6162 \$153 \$1918 \$3709 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$6163 \$153 \$153 \$3606 \$4020 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6164 \$16 \$2576 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6167 \$153 \$4080 \$4148 \$4215 \$4160 \$4110 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$6168 \$153 \$4082 \$4110 \$4215 \$4148 \$4160 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$6169 \$153 \$4148 \$4160 \$4231 \$4110 \$4215 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$6170 \$16 \$4231 \$16 \$153 \$4162 VNB sky130_fd_sc_hd__clkbuf_2
X$6172 \$16 \$4162 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6173 \$153 \$4185 \$4111 \$3572 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6174 \$16 \$3621 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6177 \$16 \$3572 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6178 \$16 \$4162 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6179 \$16 \$3811 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6180 \$153 \$4247 \$3079 \$4216 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6181 \$153 \$4086 \$4111 \$3480 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6182 \$16 \$3480 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6183 \$153 \$3877 \$4111 \$3492 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6184 \$16 \$3492 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6185 \$16 \$3386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6186 \$16 \$3492 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6189 \$153 \$4298 \$3354 \$4216 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6190 \$16 \$4229 \$4014 \$4273 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$6191 \$153 \$4248 \$3101 \$4068 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6192 \$153 \$4274 \$3954 \$3621 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6194 \$153 \$4217 \$3955 \$3492 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6196 \$153 \$4217 \$3354 \$3937 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6197 \$153 \$4218 \$3955 \$3620 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6198 \$153 \$4218 \$3645 \$3937 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6199 \$16 \$3620 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6201 \$16 \$4249 \$16 \$153 \$3783 VNB sky130_fd_sc_hd__clkbuf_2
X$6202 \$16 \$4249 \$16 \$153 \$4275 VNB sky130_fd_sc_hd__clkbuf_2
X$6203 \$153 \$4250 \$3079 \$4300 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6204 \$16 \$3621 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6206 \$16 \$3270 \$3978 \$3369 \$237 \$16 \$153 VNB sky130_fd_sc_hd__mux2_1
X$6207 \$16 \$3621 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6208 \$16 \$4249 \$16 \$153 \$4014 VNB sky130_fd_sc_hd__clkbuf_2
X$6209 \$153 \$4251 \$3354 \$4300 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6210 \$153 \$3956 \$5349 \$4043 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$6211 \$16 \$3386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6212 \$153 \$4219 \$4163 \$3386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6214 \$153 \$4219 \$3435 \$4164 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6215 \$16 \$3480 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6216 \$153 \$4220 \$4163 \$3620 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6217 \$153 \$4220 \$3645 \$4164 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6218 \$153 \$4192 \$3504 \$4164 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6219 \$153 \$4136 \$3101 \$3884 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6220 \$16 \$3620 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6223 \$153 \$4252 \$3645 \$4232 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6224 \$153 \$4137 \$3556 \$4232 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6225 \$16 \$3886 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6226 \$153 \$4221 \$4194 \$3572 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6228 \$153 \$4221 \$3101 \$4232 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6229 \$153 \$153 \$3504 \$4233 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6231 \$16 \$16 \$153 VNB sky130_fd_sc_hd__conb_1
X$6232 \$153 \$153 \$3556 \$4233 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6233 \$153 \$153 \$3645 \$4233 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6234 \$16 \$3716 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6235 \$16 \$3962 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6236 \$16 \$3335 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6237 \$153 \$3335 \$3889 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$6238 \$153 \$153 \$3919 \$4071 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6240 \$153 \$3789 \$3958 \$3731 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6241 \$153 \$153 \$3716 \$4071 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6242 \$153 \$4222 \$4254 \$3791 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6243 \$153 \$4222 \$3919 \$4234 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6244 \$16 \$3814 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6245 \$16 \$3788 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6246 \$16 \$4276 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6248 \$16 \$4093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6249 \$16 \$4093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6250 \$16 \$3852 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6251 \$153 \$4255 \$3763 \$4234 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6252 \$153 \$4277 \$4165 \$3852 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6253 \$153 \$4278 \$4165 \$3791 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6254 \$153 \$4197 \$3788 \$4235 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6256 \$153 \$3790 \$4126 \$4140 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$6257 \$16 \$3791 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6258 \$153 \$4198 \$4256 \$3791 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6259 \$16 \$4126 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6260 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$6261 \$16 \$3852 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6262 \$153 \$4279 \$4256 \$3852 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6265 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$6266 \$16 \$4415 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6267 \$16 \$3731 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6268 \$153 \$4280 \$4257 \$3731 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6269 \$153 \$4199 \$3858 \$3773 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6270 \$16 \$4258 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6271 \$16 \$4258 \$4015 \$4281 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$6272 \$153 \$3670 \$5264 \$4281 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$6273 \$16 \$3960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6276 \$153 \$4282 \$4323 \$3889 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6277 \$153 \$4282 \$3962 \$4236 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6278 \$153 \$4259 \$3651 \$4236 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6279 \$16 \$3889 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6280 \$153 \$4200 \$3962 \$3609 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6281 \$16 \$3889 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6282 \$153 \$4202 \$3939 \$4024 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6284 \$153 \$4283 \$4260 \$3889 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6285 \$16 \$3792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6286 \$16 \$4141 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6287 \$16 \$3731 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6288 \$153 \$4224 \$4260 \$3731 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6289 \$153 \$4224 \$3788 \$4237 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6290 \$153 \$4204 \$3788 \$4024 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6292 \$153 \$4261 \$3651 \$4237 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6293 \$16 \$3086 \$4262 \$3752 \$3704 \$16 \$153 VNB sky130_fd_sc_hd__mux2_1
X$6295 \$16 \$4263 \$16 \$153 \$4258 VNB sky130_fd_sc_hd__clkbuf_2
X$6296 \$16 \$4238 \$16 \$153 \$4016 VNB sky130_fd_sc_hd__clkbuf_2
X$6297 \$153 \$4238 \$4265 \$4225 \$4239 \$4266 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$6298 \$153 \$4264 \$4266 \$4225 \$4239 \$4265 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$6299 \$153 \$4239 \$4266 \$4026 \$4265 \$4225 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$6301 \$153 \$4226 \$4094 \$3721 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6302 \$153 \$4226 \$3676 \$4072 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6303 \$153 \$4240 \$4094 \$3691 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6304 \$153 \$4240 \$3142 \$4072 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6305 \$16 \$3721 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6306 \$16 \$4324 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6307 \$16 \$4093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6309 \$16 \$4093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6310 \$16 \$3826 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6311 \$153 \$4169 \$4017 \$3826 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6312 \$16 \$4139 \$16 \$153 \$3895 VNB sky130_fd_sc_hd__inv_1
X$6313 \$16 \$4139 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6315 \$16 \$4129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6316 \$153 \$4227 \$4017 \$4129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6317 \$153 \$4227 \$3986 \$3895 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6318 \$16 \$3691 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6321 \$16 \$3680 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6322 \$153 \$4284 \$4095 \$3898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6323 \$16 \$3898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6325 \$16 \$4057 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6326 \$153 \$4285 \$4095 \$4057 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6328 \$16 \$4011 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6329 \$16 \$4011 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6330 \$153 \$4061 \$3860 \$3775 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6331 \$16 \$4168 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6333 \$153 \$3829 \$4414 \$3775 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6335 \$16 \$3721 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6336 \$153 \$4286 \$4267 \$3721 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6337 \$16 \$4258 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6338 \$16 \$3680 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6339 \$153 \$4287 \$4267 \$3680 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6340 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$6341 \$16 \$3721 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6343 \$153 \$4288 \$4268 \$3721 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6344 \$16 \$4129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6345 \$153 \$4289 \$4268 \$4129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6346 \$153 \$4290 \$4268 \$3691 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6347 \$16 \$4129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6348 \$16 \$4376 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6349 \$16 \$3602 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6351 \$16 \$3680 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6353 \$153 \$4065 \$3860 \$3899 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6354 \$153 \$4291 \$4172 \$3602 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6355 \$16 \$3826 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6356 \$16 \$4092 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6358 \$16 \$3721 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6359 \$153 \$4292 \$4172 \$3721 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6360 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$6362 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$6363 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$6364 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$6365 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$6367 \$153 \$4293 \$4241 \$3766 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6368 \$16 \$3766 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6369 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$6371 \$153 \$4293 \$3478 \$4066 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6372 \$153 \$4441 \$3490 \$4066 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6373 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$6374 \$153 \$4294 \$4241 \$3571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6375 \$153 \$4294 \$3422 \$4066 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6376 \$16 \$3571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6377 \$16 \$4320 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6378 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$6380 \$153 \$4243 \$4158 \$3766 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6381 \$153 \$4326 \$4158 \$3473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6382 \$153 \$4327 \$4158 \$3385 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6383 \$16 \$4229 \$16 \$153 \$4067 VNB sky130_fd_sc_hd__inv_1
X$6384 \$16 \$4229 \$4144 \$4311 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$6386 \$153 \$4158 \$4179 \$4311 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$6387 \$153 \$4295 \$4143 \$3709 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6388 \$16 \$3709 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6390 \$153 \$4295 \$3606 \$4328 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6391 \$153 \$4270 \$3394 \$4328 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6392 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$6395 \$153 \$4159 \$4143 \$3571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6396 \$16 \$4181 \$16 \$153 \$3686 VNB sky130_fd_sc_hd__clkbuf_2
X$6397 \$153 \$4244 \$3947 \$3385 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6398 \$153 \$3947 \$5125 \$4296 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$6399 \$16 \$4106 \$4144 \$4296 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$6402 \$16 \$3766 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6404 \$153 \$3838 \$5349 \$4271 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$6405 \$16 \$4181 \$16 \$153 \$4144 VNB sky130_fd_sc_hd__clkbuf_2
X$6407 \$16 \$3616 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6408 \$153 \$4147 \$3838 \$3473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6409 \$16 \$3473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6411 \$153 \$4330 \$3389 \$4329 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6412 \$16 \$3766 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6413 \$16 \$4146 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6415 \$153 \$4297 \$4319 \$3571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6416 \$153 \$4297 \$3422 \$4230 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6417 \$16 \$3571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6418 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$6420 \$153 \$4331 \$4319 \$3709 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6421 \$16 \$3709 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6422 \$16 \$4246 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6423 \$16 \$3886 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6426 \$153 \$4332 \$3389 \$4230 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6427 \$16 \$4620 \$16 \$153 \$4020 VNB sky130_fd_sc_hd__clkbuf_2
X$6429 \$16 \$2793 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6430 \$16 \$2936 \$16 \$153 \$4078 VNB sky130_fd_sc_hd__clkbuf_2
X$6431 \$16 \$2793 \$16 \$153 \$4184 VNB sky130_fd_sc_hd__clkbuf_2
X$6432 \$16 \$2576 \$16 \$153 \$4272 VNB sky130_fd_sc_hd__clkbuf_2
X$6434 \$153 \$4333 \$4160 \$4215 \$4148 \$4110 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$6435 \$16 \$2936 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6437 \$153 \$4160 \$4110 \$4334 \$4148 \$4215 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$6438 \$16 \$4272 \$16 \$153 \$4148 VNB sky130_fd_sc_hd__clkbuf_2
X$6441 \$16 \$4333 \$16 \$153 \$3778 VNB sky130_fd_sc_hd__clkbuf_2
X$6442 \$16 \$4320 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6444 \$153 \$4335 \$4321 \$3621 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6445 \$16 \$4334 \$16 \$153 \$3879 VNB sky130_fd_sc_hd__clkbuf_2
X$6447 \$153 \$4247 \$4321 \$3573 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6448 \$16 \$3573 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6450 \$153 \$4361 \$3504 \$4216 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6452 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$6454 \$153 \$4298 \$4321 \$3492 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6455 \$153 \$4336 \$3435 \$4216 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6457 \$16 \$4229 \$16 \$153 \$4068 VNB sky130_fd_sc_hd__inv_1
X$6458 \$153 \$4248 \$3954 \$3572 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6460 \$16 \$4178 \$4014 \$4312 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$6462 \$153 \$3955 \$4269 \$4312 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$6463 \$153 \$4274 \$3608 \$4068 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6464 \$153 \$4337 \$3079 \$4338 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6465 \$16 \$3572 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6466 \$16 \$3492 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6468 \$153 \$4450 \$3435 \$4338 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6469 \$16 \$3621 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6470 \$16 \$5388 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6471 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$6472 \$16 \$4421 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6475 \$153 \$4299 \$4322 \$3621 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6476 \$153 \$4299 \$3608 \$4300 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6477 \$16 \$4421 \$16 \$153 \$4300 VNB sky130_fd_sc_hd__inv_1
X$6478 \$153 \$4313 \$4322 \$3386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6479 \$153 \$4339 \$3504 \$4300 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6480 \$16 \$3386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6482 \$153 \$4313 \$3435 \$4300 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6483 \$16 \$4249 \$16 \$153 \$3957 VNB sky130_fd_sc_hd__clkbuf_2
X$6484 \$16 \$5349 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6485 \$16 \$4106 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6486 \$16 \$3270 \$4340 \$3372 \$1099 \$16 \$153 VNB sky130_fd_sc_hd__mux2_1
X$6487 \$153 \$4453 \$3556 \$4164 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6488 \$16 \$3270 \$4668 \$3452 \$556 \$16 \$153 VNB sky130_fd_sc_hd__mux2_1
X$6490 \$16 \$3620 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6491 \$153 \$4341 \$3079 \$4363 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6494 \$153 \$4194 \$4246 \$4193 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$6495 \$153 \$4252 \$4194 \$3620 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6496 \$16 \$3886 \$16 \$153 \$4232 VNB sky130_fd_sc_hd__inv_1
X$6498 \$153 \$4116 \$3354 \$4232 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6499 \$153 \$4138 \$3504 \$4232 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6500 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$6502 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$6503 \$16 \$4620 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6504 \$153 \$4342 \$3608 \$4232 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6505 \$16 \$3572 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6506 \$16 \$4620 \$16 \$153 \$4233 VNB sky130_fd_sc_hd__clkbuf_2
X$6508 \$153 \$153 \$3079 \$4233 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6509 \$153 \$153 \$3608 \$4233 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6510 \$153 \$153 \$3101 \$4233 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6511 \$16 \$3344 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6513 \$16 \$3284 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6515 \$153 \$3284 \$4048 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$6516 \$16 \$3731 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6517 \$16 \$3792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6518 \$16 \$16 \$153 VNB sky130_fd_sc_hd__conb_1
X$6519 \$153 \$153 \$3858 \$4071 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6520 \$153 \$153 \$3763 \$4071 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6521 \$153 \$153 \$3939 \$4071 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6522 \$16 \$3791 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6524 \$153 \$4343 \$4254 \$3889 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6525 \$16 \$3889 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6526 \$16 \$3852 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6527 \$153 \$4255 \$4254 \$3852 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6528 \$153 \$4195 \$3651 \$4234 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6530 \$153 \$4314 \$3962 \$3160 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6532 \$16 \$3791 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6533 \$153 \$4277 \$3763 \$4235 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6535 \$16 \$3814 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6536 \$153 \$4301 \$4165 \$3814 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6537 \$153 \$4301 \$3651 \$4235 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6539 \$153 \$4150 \$4256 \$3960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6541 \$16 \$3731 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6542 \$153 \$4344 \$3962 \$4167 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6543 \$153 \$4302 \$4256 \$3731 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6544 \$153 \$4279 \$3763 \$4167 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6545 \$153 \$4345 \$4257 \$3814 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6546 \$16 \$3814 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6547 \$16 \$4048 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6550 \$153 \$4346 \$4257 \$4048 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6551 \$16 \$5264 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6552 \$16 \$3814 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6553 \$16 \$3889 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6554 \$16 \$3960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6555 \$153 \$4259 \$4323 \$3814 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6557 \$16 \$3731 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6558 \$16 \$3852 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6559 \$153 \$4315 \$3763 \$4236 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6561 \$153 \$4315 \$4323 \$3852 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6562 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$6563 \$16 \$4303 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6564 \$16 \$3960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6565 \$153 \$4304 \$4260 \$3960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6567 \$153 \$4304 \$3716 \$4237 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6568 \$16 \$4262 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6569 \$16 \$4203 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6570 \$16 \$4092 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6572 \$153 \$4283 \$3962 \$4237 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6574 \$16 \$4316 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6575 \$16 \$3814 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6576 \$153 \$4261 \$4260 \$3814 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6577 \$16 \$3086 \$4303 \$3528 \$245 \$16 \$153 VNB sky130_fd_sc_hd__mux2_1
X$6578 \$16 \$2793 \$16 \$153 \$4317 VNB sky130_fd_sc_hd__clkbuf_2
X$6579 \$16 \$2576 \$16 \$153 \$4305 VNB sky130_fd_sc_hd__clkbuf_2
X$6580 \$16 \$4264 \$16 \$153 \$4011 VNB sky130_fd_sc_hd__clkbuf_2
X$6581 \$16 \$4347 \$16 \$153 \$4266 VNB sky130_fd_sc_hd__clkbuf_2
X$6584 \$153 \$4263 \$4239 \$4225 \$4265 \$4266 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$6585 \$153 \$4239 \$4265 \$4348 \$4266 \$4225 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$6586 \$16 \$4225 \$4266 \$4239 \$4265 \$16 \$153 \$4349 VNB
+ sky130_fd_sc_hd__and4_2
X$6587 \$16 \$4324 \$16 \$153 \$4072 VNB sky130_fd_sc_hd__inv_1
X$6588 \$153 \$4306 \$4094 \$3898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6589 \$153 \$4306 \$3860 \$4072 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6592 \$153 \$4307 \$4094 \$3680 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6593 \$153 \$4307 \$3719 \$4072 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6594 \$16 \$4139 \$3988 \$4308 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$6595 \$16 \$4324 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6597 \$153 \$4170 \$4017 \$3680 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6598 \$16 \$3680 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6599 \$16 \$4780 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6600 \$16 \$4780 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6603 \$153 \$4309 \$4017 \$3691 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6604 \$153 \$4309 \$3142 \$3895 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6605 \$153 \$4318 \$4095 \$3680 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6606 \$153 \$4127 \$3893 \$4379 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6607 \$16 \$3691 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6608 \$16 \$4415 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6609 \$16 \$4415 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6611 \$153 \$4350 \$3719 \$4369 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6613 \$16 \$3602 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6614 \$153 \$4351 \$4325 \$3602 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6615 \$153 \$4352 \$3860 \$4369 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6617 \$16 \$4057 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6618 \$153 \$4353 \$4267 \$4057 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6621 \$16 \$3898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6622 \$153 \$4354 \$4267 \$3898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6623 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$6624 \$16 \$3602 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6625 \$153 \$4355 \$4268 \$3602 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6626 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$6628 \$16 \$4316 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6629 \$153 \$3683 \$3719 \$4171 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6632 \$16 \$3691 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6633 \$153 \$3760 \$3676 \$4171 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6634 \$153 \$3835 \$3986 \$4171 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6635 \$153 \$4310 \$4172 \$4129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6636 \$153 \$4310 \$3986 \$4173 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6637 \$153 \$4356 \$3719 \$4173 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6640 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$6641 \$16 \$3898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6642 \$153 \$4357 \$4172 \$3898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6644 \$153 \$4292 \$3676 \$4173 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6645 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$6646 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$6647 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$6648 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$6650 \$153 \$3654 \$3494 \$3709 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6652 \$153 \$3588 \$3478 \$3420 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6653 \$153 \$3654 \$3606 \$3420 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6654 \$153 \$3685 \$3389 \$3420 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6655 \$16 \$3385 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6656 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$6659 \$153 \$3626 \$3307 \$3420 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6660 \$153 \$3627 \$3490 \$3208 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6661 \$153 \$3628 \$3540 \$3208 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6663 \$153 \$3629 \$3389 \$3331 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6665 \$153 \$3424 \$3495 \$3615 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6667 \$16 \$3615 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6669 \$153 \$3655 \$3497 \$3616 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6670 \$16 \$3616 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6672 \$153 \$3630 \$3478 \$3426 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6673 \$153 \$3798 \$3606 \$3426 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6674 \$153 \$3446 \$3394 \$3426 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6675 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$6677 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$6678 \$153 \$3631 \$3389 \$3578 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6679 \$153 \$3579 \$3407 \$3766 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6680 \$153 \$3589 \$3407 \$3615 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6681 \$153 \$3589 \$3307 \$3578 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6682 \$16 \$3615 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6684 \$153 \$3656 \$3408 \$3615 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6686 \$153 \$3657 \$3499 \$3615 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6687 \$153 \$3431 \$3499 \$3385 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6688 \$16 \$3385 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6689 \$16 \$3615 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6690 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$6692 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$6693 \$153 \$3346 \$3410 \$3385 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6694 \$16 \$3385 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6696 \$16 \$2743 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6697 \$16 \$3658 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6698 \$153 \$3580 \$3410 \$3571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6699 \$153 \$3590 \$3540 \$3334 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6700 \$16 \$3571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6703 \$16 \$2743 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6704 \$153 \$3632 \$3394 \$3607 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6705 \$153 \$3303 \$1792 \$2743 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6706 \$153 \$3118 \$1547 \$2743 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6707 \$153 \$1436 \$3616 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$6708 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6709 \$16 \$1436 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6710 \$16 \$1538 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6713 \$153 \$3591 \$3659 \$3449 \$3633 \$3634 \$3618 \$3592 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$6714 \$153 \$3591 \$3619 \$3450 \$3617 \$3635 \$3516 \$3592 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$6715 \$16 \$3660 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6716 \$153 \$2991 \$1895 \$3269 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6717 \$16 \$3618 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6720 \$16 \$3636 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6721 \$16 \$3692 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6723 \$153 \$3637 \$3608 \$3336 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6724 \$16 \$3621 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6725 \$16 \$3572 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6726 \$16 \$3634 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6727 \$16 \$3638 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6728 \$153 \$3661 \$3412 \$3620 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6729 \$16 \$3692 \$16 \$153 \$3583 VNB sky130_fd_sc_hd__inv_1
X$6730 \$153 \$3639 \$3608 \$3583 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6731 \$16 \$3620 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6732 \$16 \$3692 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6733 \$16 \$3635 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6735 \$16 \$3696 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6737 \$153 \$3640 \$3645 \$3583 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6739 \$153 \$3641 \$3101 \$3583 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6740 \$153 \$3662 \$3556 \$3583 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6741 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$6742 \$153 \$3642 \$3101 \$3337 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6744 \$153 \$3643 \$3608 \$3337 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6746 \$153 \$3644 \$3645 \$3337 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6747 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$6748 \$153 \$3593 \$3413 \$3621 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6750 \$153 \$3593 \$3608 \$3339 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6752 \$153 \$3594 \$3542 \$3480 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6754 \$16 \$3480 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6755 \$16 \$3415 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6756 \$153 \$3594 \$3504 \$3506 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6757 \$153 \$3663 \$3542 \$3543 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6758 \$16 \$3572 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6759 \$153 \$3664 \$3493 \$3572 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6761 \$16 \$3572 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6762 \$16 \$3646 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6763 \$153 \$3665 \$3493 \$3480 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6764 \$153 \$3665 \$3504 \$3340 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6765 \$16 \$3480 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6766 \$153 \$3647 \$3556 \$3436 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6767 \$153 \$3401 \$3574 \$3573 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6769 \$153 \$3648 \$3608 \$3436 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6770 \$153 \$1544 \$3480 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$6771 \$16 \$16 \$153 VNB sky130_fd_sc_hd__conb_1
X$6772 \$16 \$1544 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6773 \$16 \$3335 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6774 \$153 \$1677 \$3572 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$6776 \$16 \$1677 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6777 \$16 \$1488 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6778 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6779 \$153 \$3280 \$1482 \$3645 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6780 \$153 \$3335 \$2016 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$6782 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6783 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6784 \$16 \$3272 \$3772 \$3138 \$242 \$16 \$153 VNB sky130_fd_sc_hd__mux2_1
X$6786 \$153 \$3516 \$1482 \$1558 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6787 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6788 \$153 \$3546 \$1482 \$1924 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6789 \$153 \$3223 \$1482 \$3556 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6790 \$16 \$1924 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6791 \$16 \$1878 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6792 \$16 \$2105 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6794 \$16 \$2098 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6795 \$153 \$3666 \$3281 \$1756 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6796 \$153 \$3595 \$1715 \$3341 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6797 \$16 \$3161 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6799 \$16 \$2105 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6800 \$153 \$3667 \$3211 \$2105 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6801 \$16 \$1933 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6802 \$16 \$3358 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6803 \$16 \$3210 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6804 \$16 \$2016 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6806 \$153 \$3668 \$3211 \$2016 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6807 \$16 \$3272 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6809 \$16 \$3814 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6810 \$16 \$2016 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6811 \$153 \$3669 \$3622 \$3814 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6812 \$153 \$3596 \$1715 \$3246 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6813 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$6814 \$16 \$2016 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6816 \$153 \$3597 \$3140 \$2016 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6817 \$153 \$3545 \$2438 \$3162 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6818 \$153 \$3597 \$1715 \$3162 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6819 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$6820 \$153 \$3525 \$2438 \$3317 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6821 \$153 \$3526 \$1868 \$3317 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6823 \$153 \$3671 \$3670 \$3731 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6824 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$6825 \$16 \$3731 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6826 \$153 \$3672 \$3649 \$3731 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6827 \$153 \$3650 \$3651 \$3609 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6829 \$153 \$3652 \$3788 \$3610 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6831 \$16 \$3310 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6832 \$16 \$3310 \$16 \$153 \$3530 VNB sky130_fd_sc_hd__clkbuf_2
X$6833 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6834 \$153 \$3575 \$1482 \$4414 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6835 \$16 \$3241 \$16 \$153 \$3511 VNB sky130_fd_sc_hd__clkbuf_2
X$6836 \$16 \$3241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6837 \$153 \$3530 \$3673 \$3456 \$3598 \$3653 \$3601 \$3511 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$6839 \$16 \$3576 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6840 \$16 \$3674 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6842 \$153 \$3611 \$3651 \$3610 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6843 \$16 \$3086 \$3248 \$3529 \$2546 \$16 \$153 VNB sky130_fd_sc_hd__mux2_1
X$6844 \$16 \$3688 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6845 \$16 \$3676 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6846 \$153 \$3600 \$4414 \$3461 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6847 \$153 \$3677 \$3719 \$3461 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6848 \$153 \$3675 \$1482 \$2000 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6850 \$153 \$3601 \$1482 \$2265 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6852 \$153 \$3508 \$2093 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$6853 \$153 \$3678 \$3795 \$3602 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6855 \$16 \$3587 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6857 \$153 \$3587 \$3721 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$6858 \$16 \$1860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6859 \$16 \$3691 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6860 \$153 \$3373 \$3691 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$6861 \$153 \$3188 \$1936 \$3167 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6862 \$16 \$3373 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6865 \$153 \$3600 \$3705 \$4057 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6866 \$16 \$3680 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6867 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$6868 \$153 \$3464 \$2269 \$3342 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6869 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$6870 \$153 \$3613 \$3565 \$3612 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6871 \$153 \$3465 \$2000 \$3192 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6873 \$153 \$3613 \$3623 \$3602 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6874 \$153 \$3466 \$2271 \$3192 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6876 \$153 \$3467 \$2269 \$2931 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6877 \$153 \$3681 \$3624 \$3602 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6878 \$16 \$3602 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6879 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$6881 \$16 \$1860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6882 \$153 \$3604 \$3252 \$1860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6883 \$153 \$3604 \$2000 \$3169 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6884 \$16 \$3602 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6885 \$153 \$3682 \$3722 \$3602 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6887 \$153 \$3470 \$2271 \$3328 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6889 \$153 \$3683 \$3625 \$3680 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6890 \$153 \$3614 \$3625 \$3602 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6892 \$16 \$3898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6893 \$153 \$3684 \$3625 \$3898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6894 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$6897 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$6898 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$6899 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$6900 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$6901 \$153 \$3685 \$3494 \$3616 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6902 \$16 \$3616 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6903 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$6905 \$153 \$3213 \$3708 \$3385 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6906 \$153 \$3626 \$3494 \$3615 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6907 \$16 \$3692 \$3686 \$3734 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$6908 \$16 \$3692 \$16 \$153 \$3420 VNB sky130_fd_sc_hd__inv_1
X$6909 \$153 \$3629 \$3495 \$3616 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6911 \$153 \$3723 \$3478 \$3331 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6912 \$153 \$3735 \$3495 \$3709 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6913 \$16 \$3841 \$16 \$153 \$3331 VNB sky130_fd_sc_hd__inv_1
X$6914 \$16 \$3709 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6915 \$16 \$3841 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6917 \$153 \$3630 \$3497 \$3766 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6918 \$16 \$3766 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6919 \$16 \$3709 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6921 \$16 \$3686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6923 \$153 \$3736 \$3497 \$3615 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6924 \$16 \$3615 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6926 \$153 \$3737 \$3407 \$3709 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6927 \$153 \$3631 \$3407 \$3616 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6928 \$16 \$3714 \$3686 \$3738 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$6930 \$16 \$3714 \$16 \$153 \$3578 VNB sky130_fd_sc_hd__inv_1
X$6931 \$16 \$3616 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6932 \$16 \$3714 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6934 \$153 \$3693 \$3408 \$3766 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6935 \$153 \$3693 \$3478 \$3476 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6936 \$16 \$3616 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6937 \$16 \$3766 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6939 \$153 \$3656 \$3307 \$3476 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6940 \$153 \$3657 \$3307 \$3409 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6943 \$153 \$3694 \$3499 \$3766 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6944 \$153 \$3694 \$3478 \$3409 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6945 \$16 \$3766 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6946 \$16 \$3761 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6947 \$153 \$3695 \$3410 \$3766 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6948 \$153 \$3695 \$3478 \$3334 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6952 \$16 \$3658 \$16 \$153 \$3334 VNB sky130_fd_sc_hd__inv_1
X$6953 \$16 \$3658 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6955 \$153 \$3724 \$3389 \$3334 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6956 \$153 \$3739 \$3725 \$3571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6957 \$16 \$3571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6959 \$153 \$3740 \$3725 \$3474 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6960 \$16 \$3474 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6961 \$16 \$2743 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6964 \$153 \$3741 \$3725 \$3616 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6965 \$16 \$232 \$16 \$153 \$2793 VNB sky130_fd_sc_hd__clkbuf_2
X$6966 \$16 \$232 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6967 \$153 \$3591 \$3742 \$3365 \$3710 \$3711 \$3726 \$3592 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$6968 \$16 \$3712 \$4134 \$3659 \$553 \$16 \$153 VNB sky130_fd_sc_hd__mux2_1
X$6969 \$16 \$3241 \$16 \$153 \$3592 VNB sky130_fd_sc_hd__clkbuf_2
X$6971 \$16 \$3712 \$3696 \$3619 \$208 \$16 \$153 VNB sky130_fd_sc_hd__mux2_1
X$6972 \$153 \$3637 \$3412 \$3621 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6973 \$153 \$3582 \$3412 \$3543 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6974 \$16 \$3638 \$16 \$153 \$3336 VNB sky130_fd_sc_hd__inv_1
X$6975 \$16 \$3543 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6978 \$153 \$3639 \$3713 \$3621 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6980 \$153 \$3640 \$3713 \$3620 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6981 \$153 \$3641 \$3713 \$3572 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6982 \$16 \$3620 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6983 \$16 \$3572 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6984 \$16 \$3492 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6987 \$153 \$3642 \$3502 \$3572 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6989 \$153 \$3643 \$3502 \$3621 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6990 \$16 \$3621 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6991 \$16 \$3572 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6993 \$16 \$3543 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6994 \$153 \$3697 \$3413 \$3572 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$6996 \$16 \$3621 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6997 \$16 \$3620 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$6998 \$153 \$3697 \$3101 \$3339 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$6999 \$16 \$3572 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7000 \$16 \$5183 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7001 \$153 \$3698 \$3542 \$3621 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7002 \$16 \$3714 \$16 \$153 \$3506 VNB sky130_fd_sc_hd__inv_1
X$7003 \$16 \$3621 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7005 \$153 \$3744 \$3542 \$3572 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7008 \$153 \$3727 \$3645 \$3506 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7009 \$153 \$3663 \$3556 \$3506 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7010 \$16 \$3997 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7011 \$16 \$3997 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7013 \$153 \$3664 \$3101 \$3340 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7014 \$153 \$3745 \$3493 \$3621 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7015 \$16 \$3621 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7016 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$7018 \$153 \$3647 \$3574 \$3543 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7019 \$16 \$3543 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7020 \$153 \$3728 \$3645 \$3436 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7021 \$153 \$3729 \$3079 \$3585 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7022 \$153 \$1673 \$3492 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$7024 \$16 \$1673 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7025 \$16 \$3651 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7026 \$16 \$1895 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7027 \$16 \$1954 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7028 \$153 \$3730 \$3556 \$3585 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7029 \$153 \$1488 \$3621 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$7031 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7032 \$153 \$3635 \$1482 \$3651 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7035 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7036 \$153 \$3411 \$1482 \$1613 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7038 \$153 \$3867 \$1482 \$2438 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7039 \$153 \$3726 \$1482 \$1868 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7040 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7041 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7043 \$153 \$3636 \$1482 \$1712 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7044 \$153 \$3699 \$3939 \$3160 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7045 \$153 \$3700 \$3715 \$3731 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7046 \$16 \$1756 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7047 \$16 \$3731 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7048 \$153 \$3666 \$1712 \$3341 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7049 \$16 \$3273 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7052 \$153 \$3701 \$3716 \$3160 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7053 \$153 \$3746 \$3790 \$3731 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7054 \$153 \$3667 \$2438 \$3203 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7055 \$153 \$3668 \$1715 \$3203 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7057 \$16 \$3852 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7058 \$153 \$3669 \$3651 \$3732 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7060 \$153 \$3702 \$3622 \$3852 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7061 \$153 \$3702 \$3763 \$3732 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7062 \$153 \$3819 \$3939 \$3732 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7063 \$153 \$3747 \$3717 \$3814 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7064 \$16 \$3814 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7066 \$16 \$3852 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7068 \$153 \$3748 \$3717 \$3852 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7070 \$16 \$3852 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7071 \$153 \$3749 \$3670 \$3852 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7072 \$153 \$3563 \$1715 \$3317 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7073 \$153 \$3749 \$3763 \$3891 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7075 \$16 \$3852 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7077 \$153 \$3750 \$3649 \$3852 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7079 \$16 \$3852 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7080 \$153 \$3751 \$3718 \$3852 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7081 \$153 \$3652 \$3718 \$3731 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7082 \$16 \$3418 \$16 \$153 \$3086 VNB sky130_fd_sc_hd__clkbuf_2
X$7085 \$153 \$3733 \$3962 \$3610 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7087 \$153 \$3530 \$3752 \$3559 \$3599 \$3689 \$3533 \$3511 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$7088 \$153 \$3530 \$3753 \$3688 \$3674 \$3703 \$3566 \$3511 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$7089 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7090 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7093 \$153 \$3703 \$1482 \$3676 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7094 \$153 \$3754 \$1482 \$3719 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7095 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7097 \$153 \$3199 \$4057 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$7099 \$153 \$3824 \$3676 \$3586 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7100 \$153 \$3720 \$1860 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$7101 \$153 \$3678 \$3565 \$3586 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7102 \$16 \$3720 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7103 \$153 \$3165 \$3705 \$3691 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7105 \$153 \$3379 \$2271 \$3167 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7106 \$16 \$3720 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7108 \$153 \$3677 \$3705 \$3680 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7109 \$153 \$3463 \$2000 \$3342 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7111 \$153 \$3755 \$3796 \$3680 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7114 \$16 \$3691 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7115 \$153 \$3756 \$3796 \$3691 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7116 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$7117 \$16 \$3721 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7118 \$153 \$3757 \$3623 \$3721 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7119 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$7121 \$153 \$3603 \$2000 \$2931 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7124 \$16 \$3721 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7126 \$16 \$3691 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7127 \$153 \$3690 \$3624 \$3691 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7128 \$153 \$3706 \$3624 \$4057 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7129 \$153 \$3758 \$3722 \$4057 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7130 \$16 \$3691 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7132 \$153 \$3707 \$3722 \$3691 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7133 \$153 \$3707 \$3142 \$3764 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7134 \$16 \$3691 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7135 \$153 \$3759 \$3625 \$3691 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7136 \$16 \$3602 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7137 \$153 \$3605 \$2000 \$3328 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7140 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$7141 \$16 \$3721 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7142 \$153 \$3760 \$3625 \$3721 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7143 \$153 \$3383 \$2086 \$3328 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7144 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$7145 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$7146 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$7147 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$7149 \$153 \$9734 \$9875 \$9129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7151 \$153 \$9876 \$8912 \$9728 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7152 \$153 \$9877 \$8194 \$9728 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7153 \$153 \$9878 \$8885 \$9728 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7154 \$16 \$8114 \$9547 \$9894 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$7156 \$16 \$8724 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7157 \$153 \$9895 \$9831 \$8950 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7158 \$16 \$8950 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7160 \$153 \$9800 \$9831 \$9129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7161 \$153 \$9716 \$9831 \$8724 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7162 \$16 \$9129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7165 \$153 \$9448 \$9832 \$8724 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7166 \$16 \$9129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7167 \$153 \$9833 \$9543 \$8950 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7168 \$153 \$9864 \$9879 \$8724 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7169 \$16 \$8271 \$9547 \$9896 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$7172 \$153 \$9864 \$8457 \$9865 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7173 \$16 \$8724 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7174 \$153 \$9834 \$9765 \$8950 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7176 \$153 \$9834 \$8912 \$9740 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7177 \$16 \$8436 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7179 \$153 \$9897 \$9793 \$9129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7181 \$16 \$9129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7182 \$16 \$8724 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7184 \$16 \$8118 \$16 \$153 \$9866 VNB sky130_fd_sc_hd__inv_1
X$7185 \$153 \$9898 \$9793 \$8436 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7186 \$16 \$8950 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7187 \$16 \$8436 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7188 \$153 \$9835 \$9880 \$8950 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7189 \$153 \$9835 \$8912 \$9836 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7190 \$16 \$8950 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7193 \$153 \$10013 \$9880 \$9129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7194 \$16 \$8125 \$9260 \$9837 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$7195 \$153 \$9805 \$9838 \$9129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7197 \$16 \$8436 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7198 \$153 \$9806 \$9838 \$8724 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7200 \$16 \$8125 \$16 \$153 \$9867 VNB sky130_fd_sc_hd__inv_1
X$7201 \$153 \$9881 \$8912 \$9867 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7202 \$153 \$10042 \$9129 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$7203 \$153 \$9869 \$8724 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$7204 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7205 \$16 \$9869 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7207 \$153 \$9899 \$9787 \$8816 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7208 \$16 \$8816 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7209 \$153 \$9900 \$8193 \$9923 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$7210 \$16 \$9371 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7211 \$16 \$9371 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7212 \$16 \$8193 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7213 \$153 \$9901 \$9787 \$8898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7214 \$16 \$8898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7216 \$153 \$9613 \$9787 \$8556 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7217 \$153 \$9882 \$8818 \$9868 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7218 \$16 \$8139 \$16 \$153 \$9902 VNB sky130_fd_sc_hd__inv_1
X$7219 \$153 \$9839 \$9794 \$8647 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7220 \$153 \$9839 \$8614 \$9902 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7221 \$16 \$8647 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7225 \$153 \$9840 \$9795 \$8647 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7226 \$153 \$9796 \$8503 \$9883 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$7227 \$16 \$8647 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7228 \$153 \$9841 \$9796 \$8647 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7229 \$16 \$8423 \$16 \$153 \$9842 VNB sky130_fd_sc_hd__inv_1
X$7230 \$16 \$8647 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7231 \$16 \$8423 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7233 \$153 \$9841 \$8614 \$9842 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7234 \$16 \$8177 \$9400 \$9810 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$7236 \$153 \$9903 \$9811 \$8647 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7237 \$153 \$9903 \$8614 \$9586 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7238 \$153 \$9814 \$9884 \$8556 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7240 \$16 \$8556 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7241 \$16 \$9885 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7242 \$16 \$9886 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7243 \$16 \$8118 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7244 \$153 \$9843 \$9884 \$8647 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7245 \$153 \$9843 \$8614 \$9815 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7246 \$16 \$8125 \$16 \$153 \$9815 VNB sky130_fd_sc_hd__inv_1
X$7247 \$16 \$8118 \$16 \$153 \$9845 VNB sky130_fd_sc_hd__inv_1
X$7248 \$153 \$9817 \$9846 \$8728 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7251 \$153 \$9904 \$9846 \$8890 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7252 \$153 \$9847 \$8727 \$9452 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7253 \$16 \$8886 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7254 \$153 \$9905 \$9660 \$8816 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7256 \$16 \$8898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7257 \$153 \$9516 \$8610 \$9300 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7260 \$153 \$9906 \$9660 \$8898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7262 \$153 \$8364 \$9031 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$7263 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7265 \$153 \$9623 \$9732 \$9031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7267 \$16 \$8516 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7268 \$16 \$9845 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7269 \$153 \$9691 \$9732 \$9045 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7270 \$153 \$9907 \$8277 \$9746 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7272 \$153 \$153 \$9278 \$9625 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7273 \$153 \$153 \$9252 \$9625 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7275 \$16 \$8187 \$9518 \$9849 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$7276 \$16 \$8807 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7278 \$153 \$9850 \$9693 \$9253 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7279 \$153 \$9908 \$9047 \$9453 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7280 \$16 \$9275 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7281 \$153 \$9749 \$9693 \$9275 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7282 \$153 \$9870 \$8676 \$9871 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7283 \$16 \$8187 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7284 \$16 \$9031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7286 \$153 \$9851 \$9674 \$9031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7287 \$153 \$9887 \$9047 \$9695 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7289 \$153 \$9888 \$9278 \$9695 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7290 \$153 \$9818 \$9544 \$9214 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7291 \$16 \$8626 \$9518 \$9909 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$7293 \$153 \$9751 \$9544 \$9253 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7295 \$16 \$9275 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7296 \$153 \$9853 \$9752 \$9275 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7297 \$153 \$9753 \$9752 \$9214 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7298 \$16 \$8624 \$9733 \$9854 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$7300 \$16 \$9045 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7301 \$153 \$9757 \$9752 \$9045 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7302 \$16 \$8624 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7303 \$153 \$9574 \$8917 \$9521 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7304 \$153 \$9819 \$9252 \$9642 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7305 \$16 \$8807 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7306 \$153 \$9756 \$9755 \$8807 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7308 \$16 \$9031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7310 \$153 \$9889 \$9047 \$9725 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7311 \$16 \$9045 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7312 \$153 \$9855 \$9755 \$9045 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7313 \$153 \$9890 \$9174 \$9872 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7314 \$153 \$9891 \$8676 \$9872 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7315 \$16 \$8704 \$9733 \$9911 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$7317 \$16 \$9045 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7319 \$153 \$9822 \$9758 \$9188 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7320 \$153 \$9892 \$9047 \$9823 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7322 \$153 \$9912 \$9758 \$9031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7323 \$153 \$9790 \$9278 \$9823 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7324 \$16 \$8165 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7326 \$16 \$8673 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7328 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7329 \$153 \$9856 \$8340 \$8996 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7330 \$153 \$9913 \$8719 \$9873 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$7331 \$16 \$8673 \$9675 \$9873 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$7333 \$153 \$9857 \$9702 \$8927 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7334 \$16 \$8893 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7336 \$153 \$9779 \$9122 \$9759 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7337 \$153 \$9893 \$8923 \$9981 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7338 \$153 \$9914 \$9702 \$8893 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7339 \$16 \$8893 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7340 \$16 \$8927 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7342 \$153 \$9825 \$9103 \$9759 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7343 \$16 \$7996 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7344 \$16 \$8313 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7346 \$16 \$9034 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7348 \$153 \$9633 \$9676 \$8879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7349 \$153 \$9827 \$9676 \$9154 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7350 \$16 \$9154 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7351 \$16 \$8879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7352 \$16 \$8893 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7353 \$16 \$8893 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7354 \$153 \$9874 \$9677 \$8893 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7357 \$153 \$9874 \$8996 \$9592 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7359 \$16 \$9154 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7360 \$153 \$9858 \$9677 \$8879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7361 \$153 \$9858 \$8923 \$9592 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7362 \$16 \$8879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7363 \$153 \$9915 \$9726 \$9134 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7366 \$153 \$9859 \$8977 \$9708 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7368 \$16 \$8879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7369 \$153 \$9916 \$9726 \$8879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7370 \$153 \$9861 \$9726 \$9034 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7371 \$153 \$9861 \$9059 \$9708 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7372 \$16 \$9034 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7374 \$153 \$9917 \$9678 \$9034 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7375 \$153 \$9918 \$9256 \$9961 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7376 \$153 \$9919 \$9678 \$9154 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7378 \$16 \$8428 \$9562 \$9920 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$7379 \$153 \$8480 \$7180 \$8266 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7381 \$16 \$8428 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7382 \$16 \$8893 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7383 \$153 \$9921 \$9792 \$8893 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7384 \$153 \$8776 \$7375 \$8777 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7385 \$16 \$8265 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7386 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$7387 \$16 \$9034 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7388 \$153 \$9922 \$9792 \$9034 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7389 \$16 \$9035 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7392 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$7393 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$7394 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$7395 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$7396 \$153 \$9876 \$9875 \$8950 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7397 \$16 \$8950 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7398 \$16 \$8580 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7401 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$7402 \$153 \$9737 \$9875 \$8724 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7403 \$153 \$9875 \$8193 \$9894 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$7404 \$16 \$8139 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7405 \$16 \$8193 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7406 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$7407 \$153 \$9895 \$8912 \$9729 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7410 \$153 \$9945 \$8726 \$9729 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7411 \$16 \$8139 \$16 \$153 \$9729 VNB sky130_fd_sc_hd__inv_1
X$7412 \$153 \$9962 \$9832 \$8950 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7413 \$16 \$8950 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7415 \$153 \$9738 \$9832 \$9129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7416 \$153 \$9928 \$8737 \$9865 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7418 \$153 \$9928 \$9879 \$9129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7419 \$16 \$9129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7421 \$153 \$9963 \$9879 \$8950 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7422 \$16 \$8271 \$16 \$153 \$9865 VNB sky130_fd_sc_hd__inv_1
X$7423 \$16 \$8950 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7424 \$153 \$9929 \$9765 \$8436 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7426 \$16 \$8950 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7427 \$153 \$9929 \$8209 \$9740 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7428 \$153 \$9766 \$8457 \$9740 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7429 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$7430 \$16 \$8580 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7431 \$153 \$9964 \$9793 \$8950 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7432 \$153 \$9793 \$8025 \$9803 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$7434 \$153 \$9965 \$9880 \$8580 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7435 \$153 \$9966 \$9880 \$9026 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7436 \$153 \$9654 \$9880 \$8724 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7437 \$16 \$8177 \$16 \$153 \$9836 VNB sky130_fd_sc_hd__inv_1
X$7438 \$16 \$9026 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7439 \$16 \$9129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7442 \$153 \$9946 \$8209 \$9836 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7443 \$153 \$10058 \$8885 \$9867 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7444 \$153 \$9881 \$9838 \$8950 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7445 \$153 \$9339 \$8950 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$7446 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7448 \$153 \$9967 \$8340 \$8209 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7449 \$153 \$9947 \$8340 \$8737 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7450 \$153 \$9968 \$9787 \$8890 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7451 \$16 \$8114 \$9371 \$9923 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$7452 \$16 \$8890 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7455 \$153 \$9899 \$8804 \$9451 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7457 \$153 \$9901 \$8789 \$9451 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7458 \$153 \$9461 \$9787 \$8728 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7459 \$153 \$9948 \$8651 \$9868 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7460 \$153 \$9949 \$8610 \$9868 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7461 \$16 \$8556 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7465 \$153 \$9930 \$9794 \$8886 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7467 \$153 \$9795 \$8335 \$9772 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$7469 \$153 \$9931 \$9795 \$8556 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7470 \$16 \$8423 \$9371 \$9883 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$7471 \$16 \$8556 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7473 \$153 \$9931 \$8610 \$9720 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7474 \$16 \$9371 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7476 \$153 \$9932 \$9796 \$8556 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7477 \$153 \$9932 \$8610 \$9842 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7478 \$16 \$8556 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7480 \$153 \$9744 \$9811 \$8886 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7482 \$153 \$9809 \$8818 \$9842 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7483 \$16 \$8647 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7484 \$16 \$8886 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7486 \$153 \$9924 \$9884 \$8686 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7487 \$16 \$8686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7488 \$16 \$8886 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7490 \$153 \$9789 \$9884 \$8728 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7491 \$16 \$8118 \$9400 \$9844 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$7493 \$16 \$8647 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7494 \$16 \$8728 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7496 \$153 \$9925 \$9846 \$8647 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7497 \$153 \$9773 \$8614 \$9488 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7498 \$16 \$8647 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7499 \$16 \$8728 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7500 \$153 \$9969 \$9846 \$8556 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7501 \$16 \$8556 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7502 \$16 \$8890 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7506 \$16 \$8890 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7507 \$153 \$9905 \$8804 \$9746 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7508 \$153 \$6893 \$8671 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$7509 \$153 \$9907 \$9660 \$8890 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7510 \$16 \$6893 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7511 \$16 \$8364 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7512 \$16 \$10238 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7513 \$16 \$8671 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7515 \$153 \$8671 \$8807 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$7516 \$153 \$9971 \$9732 \$9253 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7518 \$153 \$9950 \$9732 \$9188 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7519 \$16 \$9188 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7522 \$153 \$9972 \$9732 \$9275 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7523 \$16 \$8187 \$16 \$153 \$9453 VNB sky130_fd_sc_hd__inv_1
X$7524 \$16 \$8673 \$9518 \$9973 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$7525 \$153 \$9926 \$9693 \$9188 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7526 \$153 \$9694 \$9693 \$9214 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7528 \$153 \$9944 \$8676 \$10216 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7529 \$153 \$9951 \$9174 \$9871 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7531 \$16 \$9253 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7532 \$153 \$9933 \$9674 \$9253 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7533 \$153 \$9933 \$9252 \$9695 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7535 \$153 \$9952 \$8676 \$9953 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7537 \$16 \$9275 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7538 \$16 \$8731 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7539 \$153 \$9934 \$8731 \$9909 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$7541 \$16 \$8807 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7542 \$153 \$9910 \$9934 \$8807 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7543 \$16 \$9275 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7545 \$153 \$9954 \$9133 \$9927 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7546 \$16 \$8626 \$16 \$153 \$9927 VNB sky130_fd_sc_hd__inv_1
X$7547 \$16 \$9253 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7548 \$16 \$8626 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7550 \$153 \$9910 \$8676 \$9927 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7551 \$16 \$9214 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7552 \$16 \$9188 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7553 \$153 \$9974 \$9752 \$9188 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7555 \$16 \$8807 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7556 \$153 \$9975 \$9752 \$8807 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7558 \$16 \$8428 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7559 \$16 \$8428 \$9733 \$9935 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$7561 \$153 \$10024 \$8666 \$9935 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$7562 \$16 \$9214 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7563 \$153 \$9976 \$9755 \$9253 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7564 \$16 \$9253 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7565 \$16 \$9642 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7566 \$16 \$9642 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7567 \$16 \$9275 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7568 \$153 \$9936 \$9755 \$9275 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7570 \$153 \$9936 \$9278 \$9725 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7572 \$16 \$8165 \$9733 \$9977 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$7573 \$153 \$9937 \$9133 \$9872 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7574 \$153 \$9938 \$9758 \$9253 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7575 \$153 \$9938 \$9252 \$9823 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7576 \$16 \$8165 \$16 \$153 \$9955 VNB sky130_fd_sc_hd__inv_1
X$7577 \$16 \$8936 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7578 \$16 \$8936 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7580 \$153 \$9978 \$9758 \$8936 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7581 \$153 \$9939 \$8842 \$9955 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7582 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7583 \$153 \$9979 \$8340 \$8965 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7584 \$153 \$9912 \$9133 \$9823 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7585 \$16 \$8965 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7586 \$16 \$8923 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7588 \$153 \$9980 \$9913 \$9035 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7589 \$16 \$8673 \$16 \$153 \$9981 VNB sky130_fd_sc_hd__inv_1
X$7590 \$16 \$8313 \$9675 \$9956 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$7591 \$153 \$9982 \$9913 \$8844 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7592 \$153 \$9940 \$8820 \$9956 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$7593 \$16 \$8844 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7595 \$153 \$9983 \$9940 \$8927 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7596 \$16 \$8893 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7597 \$16 \$7996 \$9675 \$9984 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$7598 \$153 \$9985 \$9940 \$8844 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7600 \$153 \$9561 \$9676 \$9034 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7602 \$16 \$8844 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7603 \$153 \$10085 \$8731 \$9986 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$7604 \$153 \$10130 \$9103 \$10011 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7605 \$16 \$7996 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7607 \$153 \$9957 \$8996 \$10011 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7608 \$153 \$9958 \$9256 \$10011 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7610 \$153 \$9798 \$7462 \$8429 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7612 \$153 \$9959 \$8965 \$10110 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7613 \$16 \$9154 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7614 \$16 \$8624 \$9562 \$9987 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$7615 \$153 \$9941 \$9726 \$9154 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7616 \$153 \$9941 \$9103 \$9708 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7617 \$16 \$8624 \$16 \$153 \$9988 VNB sky130_fd_sc_hd__inv_1
X$7618 \$16 \$8624 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7620 \$153 \$9706 \$9256 \$9708 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7622 \$153 \$9916 \$8923 \$9708 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7623 \$153 \$9942 \$9860 \$8893 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7624 \$16 \$8453 \$16 \$153 \$9961 VNB sky130_fd_sc_hd__inv_1
X$7625 \$16 \$8927 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7627 \$153 \$9960 \$8965 \$9961 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7628 \$153 \$9942 \$8996 \$9961 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7629 \$16 \$8704 \$9562 \$9989 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$7630 \$16 \$9154 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7632 \$153 \$9990 \$9678 \$8879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7634 \$153 \$9991 \$8666 \$9920 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$7636 \$16 \$8927 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7637 \$153 \$9943 \$9792 \$8927 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7638 \$16 \$8266 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7639 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$7641 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$7643 \$16 \$9154 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7644 \$153 \$9992 \$9792 \$9154 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7645 \$153 \$8631 \$7376 \$8777 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7647 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$7648 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$7649 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$7650 \$153 \$9283 \$9193 \$8715 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7652 \$153 \$9283 \$8638 \$9025 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7653 \$153 \$9352 \$9193 \$8828 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7654 \$16 \$8828 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7655 \$16 \$8724 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7656 \$16 \$8436 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7657 \$16 \$9026 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7659 \$153 \$9267 \$9193 \$8436 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7661 \$153 \$9330 \$8737 \$9270 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7662 \$153 \$9197 \$9196 \$8715 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7663 \$153 \$9331 \$8209 \$9270 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7664 \$16 \$8950 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7666 \$16 \$8724 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7668 \$153 \$9038 \$9196 \$9026 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7670 \$16 \$8715 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7671 \$153 \$9285 \$9130 \$8715 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7673 \$153 \$9285 \$8638 \$9136 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7674 \$153 \$9332 \$8912 \$9136 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7675 \$16 \$8950 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7678 \$153 \$9158 \$8209 \$9136 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7679 \$153 \$9353 \$9131 \$8828 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7680 \$153 \$9286 \$8457 \$9136 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7681 \$16 \$8828 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7683 \$16 \$8724 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7684 \$153 \$9288 \$9131 \$8580 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7686 \$153 \$9288 \$8194 \$9027 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7687 \$153 \$9354 \$8726 \$9321 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7689 \$153 \$9333 \$8209 \$9322 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7690 \$153 \$9323 \$9334 \$9026 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7691 \$153 \$9323 \$8726 \$9322 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7693 \$16 \$8715 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7695 \$153 \$9355 \$9334 \$8715 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7696 \$153 \$9289 \$8457 \$9029 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7698 \$153 \$9291 \$9160 \$8828 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7699 \$16 \$8436 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7700 \$153 \$9291 \$8885 \$9072 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7701 \$16 \$6903 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7704 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$7705 \$153 \$9292 \$9160 \$9129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7706 \$153 \$9292 \$8737 \$9072 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7708 \$16 \$7381 \$8635 \$9335 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$7709 \$153 \$9356 \$7547 \$9335 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$7710 \$16 \$8635 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7713 \$153 \$9203 \$9202 \$8886 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7714 \$16 \$8816 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7715 \$153 \$9204 \$9202 \$8647 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7716 \$16 \$8647 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7717 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$7718 \$153 \$9357 \$9202 \$8556 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7720 \$153 \$9293 \$8789 \$9185 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7721 \$16 \$8556 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7722 \$16 \$8556 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7723 \$16 \$8438 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7724 \$16 \$8003 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7725 \$153 \$9272 \$9001 \$8728 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7726 \$16 \$8728 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7727 \$16 \$8890 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7729 \$16 \$8886 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7730 \$153 \$9274 \$9001 \$8886 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7732 \$153 \$9337 \$8818 \$9186 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7733 \$153 \$9294 \$8789 \$8887 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7735 \$153 \$9208 \$9132 \$8816 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7736 \$153 \$9295 \$9132 \$8647 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7737 \$16 \$8647 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7738 \$16 \$8886 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7741 \$153 \$9295 \$8614 \$9111 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7742 \$153 \$9358 \$9076 \$8647 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7743 \$153 \$9359 \$9076 \$8816 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7744 \$153 \$9359 \$8804 \$9144 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7745 \$16 \$8816 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7746 \$16 \$7973 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7749 \$153 \$9338 \$8277 \$9144 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7750 \$16 \$8728 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7751 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$7753 \$153 \$9209 \$9077 \$8816 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7754 \$16 \$8816 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7755 \$16 \$8886 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7757 \$16 \$8728 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7758 \$153 \$9298 \$9077 \$8728 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7760 \$153 \$9298 \$8818 \$9146 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7762 \$153 \$9210 \$9044 \$8647 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7763 \$16 \$8647 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7764 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$7765 \$153 \$9212 \$9044 \$8816 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7766 \$153 \$9299 \$8789 \$8989 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7768 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$7770 \$153 \$153 \$8277 \$9010 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7771 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7772 \$16 \$7215 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7773 \$16 \$9339 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7774 \$153 \$9339 \$7387 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$7776 \$16 \$8126 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7777 \$16 \$8126 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7778 \$153 \$9340 \$9278 \$8126 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7780 \$16 \$8126 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7781 \$16 \$8126 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7783 \$16 \$9253 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7784 \$153 \$9341 \$8676 \$9324 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7785 \$153 \$9342 \$9174 \$9324 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7786 \$153 \$9343 \$8842 \$9324 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7787 \$153 \$9261 \$8935 \$9253 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7788 \$16 \$9253 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7789 \$16 \$7344 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7790 \$16 \$7344 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7792 \$16 \$7709 \$8819 \$9344 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$7793 \$153 \$9405 \$7903 \$9344 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$7794 \$153 \$9360 \$8900 \$9275 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7795 \$153 \$9262 \$8900 \$9253 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7797 \$16 \$8819 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7798 \$16 \$9275 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7800 \$153 \$9493 \$8917 \$8891 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7801 \$16 \$9214 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7802 \$153 \$9301 \$9081 \$9275 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7803 \$153 \$9301 \$9278 \$9276 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7804 \$16 \$7667 \$16 \$153 \$9276 VNB sky130_fd_sc_hd__inv_1
X$7806 \$153 \$9302 \$8937 \$9275 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7808 \$153 \$9302 \$9278 \$8843 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7809 \$16 \$9275 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7810 \$16 \$7495 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7811 \$16 \$9253 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7812 \$153 \$9304 \$9050 \$9253 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7813 \$153 \$9724 \$8917 \$9325 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7814 \$153 \$9304 \$9252 \$8993 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7816 \$16 \$9455 \$16 \$153 \$8960 VNB sky130_fd_sc_hd__clkbuf_2
X$7817 \$16 \$9275 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7819 \$153 \$9345 \$8842 \$9325 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7820 \$16 \$7952 \$16 \$153 \$9325 VNB sky130_fd_sc_hd__inv_1
X$7822 \$153 \$9326 \$9052 \$9275 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7824 \$16 \$9188 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7825 \$153 \$9361 \$9052 \$9188 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7826 \$16 \$7952 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7827 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$7830 \$16 \$9253 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7831 \$153 \$9308 \$9053 \$9253 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7832 \$153 \$9307 \$9278 \$8920 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7833 \$153 \$9308 \$9252 \$8920 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7834 \$153 \$9346 \$8917 \$8920 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7835 \$153 \$9327 \$8917 \$9328 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7837 \$153 \$9348 \$9347 \$9045 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7838 \$153 \$9348 \$9174 \$9328 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7840 \$16 \$8807 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7841 \$153 \$9362 \$9347 \$8807 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7842 \$153 \$9177 \$9133 \$9151 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7843 \$16 \$9275 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7846 \$16 \$7852 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7848 \$153 \$9349 \$8996 \$9152 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7849 \$153 \$9349 \$9179 \$8893 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7850 \$16 \$7386 \$16 \$153 \$9152 VNB sky130_fd_sc_hd__inv_1
X$7851 \$16 \$8893 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7852 \$16 \$7484 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7853 \$153 \$9310 \$8977 \$9152 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7855 \$16 \$9035 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7856 \$153 \$9311 \$9103 \$9152 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7859 \$153 \$9350 \$9059 \$9439 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7860 \$16 \$7709 \$8824 \$9388 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$7862 \$153 \$9351 \$9059 \$9329 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7863 \$153 \$9363 \$9441 \$8879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7864 \$153 \$9235 \$9122 \$8906 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7865 \$16 \$8879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7866 \$16 \$9034 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7867 \$16 \$9134 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7869 \$153 \$9312 \$9279 \$8893 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7870 \$153 \$9312 \$8996 \$9264 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7872 \$16 \$9154 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7873 \$153 \$9313 \$9279 \$9154 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7874 \$153 \$9313 \$9103 \$9264 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7876 \$16 \$9035 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7878 \$153 \$9314 \$9279 \$9035 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7879 \$153 \$9314 \$8977 \$9264 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7880 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$7881 \$16 \$9134 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7882 \$153 \$8845 \$8926 \$9134 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7883 \$153 \$9315 \$9059 \$8846 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7886 \$16 \$9034 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7887 \$153 \$9365 \$9364 \$9034 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7888 \$16 \$7693 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7889 \$16 \$7691 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7890 \$16 \$9035 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7891 \$153 \$9265 \$9364 \$9035 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7892 \$16 \$8844 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7893 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$7894 \$153 \$9380 \$9256 \$9239 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7896 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$7897 \$16 \$8879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7898 \$153 \$9317 \$9316 \$8879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7899 \$153 \$9317 \$8923 \$9239 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7900 \$16 \$8893 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7901 \$153 \$9218 \$9240 \$8893 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7902 \$16 \$7431 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7903 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$7905 \$153 \$9318 \$8923 \$9192 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7906 \$16 \$7695 \$16 \$153 \$9366 VNB sky130_fd_sc_hd__inv_1
X$7907 \$16 \$7695 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7909 \$153 \$9319 \$9122 \$9192 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7911 \$16 \$8844 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7912 \$16 \$9154 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7913 \$153 \$9367 \$9240 \$8844 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7915 \$153 \$9320 \$9103 \$9192 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7917 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$7918 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$7919 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$7920 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$7922 \$153 \$9194 \$9193 \$8580 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7923 \$16 \$8715 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7924 \$16 \$8580 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7927 \$153 \$9382 \$8737 \$9392 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7928 \$16 \$9129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7930 \$153 \$9266 \$9193 \$9026 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7931 \$153 \$9352 \$8885 \$9025 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7932 \$16 \$7381 \$8577 \$9383 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$7933 \$153 \$9458 \$7547 \$9383 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$7935 \$153 \$9368 \$9196 \$8950 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7936 \$153 \$8969 \$9196 \$8724 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7937 \$153 \$9393 \$8638 \$9270 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7938 \$153 \$9394 \$8726 \$9270 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7939 \$16 \$9026 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7940 \$16 \$8438 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7941 \$16 \$8003 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7943 \$153 \$9332 \$9130 \$8950 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7944 \$153 \$9412 \$9130 \$9129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7945 \$16 \$9129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7946 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$7947 \$153 \$9271 \$9131 \$9026 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7949 \$16 \$8950 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7951 \$153 \$9353 \$8885 \$9027 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7953 \$153 \$9369 \$9131 \$8724 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7954 \$153 \$9369 \$8457 \$9027 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7955 \$153 \$9475 \$8885 \$9321 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7956 \$153 \$9413 \$8737 \$9321 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7957 \$16 \$9414 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7960 \$153 \$9333 \$9334 \$8436 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7961 \$153 \$9395 \$8194 \$9322 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7962 \$16 \$8436 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7963 \$153 \$9415 \$9334 \$8724 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7964 \$153 \$9355 \$8638 \$9322 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7965 \$16 \$8828 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7966 \$16 \$8724 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7968 \$153 \$9384 \$6903 \$9290 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$7970 \$153 \$9370 \$9384 \$8436 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7971 \$153 \$9370 \$8209 \$9396 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7973 \$16 \$7381 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7974 \$16 \$7547 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7975 \$16 \$9129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7976 \$153 \$9397 \$8457 \$9396 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7978 \$153 \$9223 \$8457 \$9072 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7979 \$153 \$9398 \$8737 \$9396 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7980 \$16 \$6753 \$16 \$153 \$9396 VNB sky130_fd_sc_hd__inv_1
X$7981 \$16 \$7922 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7982 \$16 \$8635 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7983 \$153 \$9416 \$9356 \$8890 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7985 \$153 \$9224 \$8277 \$9185 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7986 \$16 \$7381 \$16 \$153 \$9417 VNB sky130_fd_sc_hd__inv_1
X$7987 \$16 \$8886 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7989 \$16 \$8890 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7990 \$16 \$7381 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7991 \$16 \$6753 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$7993 \$153 \$9385 \$8610 \$9417 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7994 \$153 \$9385 \$9356 \$8556 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$7995 \$153 \$9357 \$8610 \$9185 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7996 \$153 \$9418 \$8651 \$9417 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$7997 \$16 \$8003 \$9371 \$9419 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$7999 \$16 \$8728 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8000 \$16 \$9371 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8001 \$16 \$9371 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8002 \$16 \$8003 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8003 \$153 \$9482 \$8610 \$9186 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8004 \$153 \$9372 \$9481 \$8686 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8005 \$153 \$9372 \$8651 \$9186 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8006 \$16 \$9273 \$16 \$153 \$9371 VNB sky130_fd_sc_hd__clkbuf_2
X$8008 \$153 \$9399 \$8277 \$9373 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8010 \$153 \$9485 \$8614 \$9373 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8011 \$16 \$8816 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8012 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$8013 \$153 \$9374 \$9132 \$8890 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8014 \$153 \$9386 \$8610 \$9373 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8015 \$153 \$9296 \$8610 \$9111 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8016 \$16 \$8890 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8018 \$16 \$8556 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8019 \$16 \$8647 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8022 \$153 \$9358 \$8614 \$9144 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8023 \$16 \$7992 \$9400 \$9420 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$8024 \$153 \$9338 \$9076 \$8890 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8025 \$16 \$8890 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8026 \$16 \$7992 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8027 \$16 \$7992 \$16 \$153 \$9421 VNB sky130_fd_sc_hd__inv_1
X$8028 \$153 \$9401 \$8804 \$9421 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8030 \$153 \$9402 \$8727 \$9421 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8032 \$153 \$9297 \$8727 \$9146 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8033 \$16 \$7663 \$9400 \$9422 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$8034 \$16 \$7663 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8036 \$153 \$9423 \$9403 \$8556 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8037 \$153 \$9424 \$6903 \$9489 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$8038 \$153 \$9226 \$8277 \$8989 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8041 \$153 \$9425 \$9424 \$8816 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8042 \$16 \$6753 \$16 \$153 \$9300 VNB sky130_fd_sc_hd__inv_1
X$8043 \$16 \$8816 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8044 \$16 \$8898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8045 \$153 \$9426 \$9424 \$8898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8046 \$153 \$9336 \$8340 \$7490 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8049 \$153 \$8590 \$9404 \$8807 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8050 \$153 \$9147 \$9404 \$9253 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8052 \$153 \$9046 \$9404 \$9214 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8053 \$16 \$7793 \$8819 \$9427 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$8056 \$16 \$7793 \$16 \$153 \$8126 VNB sky130_fd_sc_hd__inv_1
X$8057 \$16 \$9214 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8058 \$16 \$9214 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8059 \$153 \$9428 \$9405 \$9214 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8060 \$153 \$9229 \$8917 \$8958 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8062 \$16 \$8819 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8063 \$16 \$7709 \$16 \$153 \$9324 VNB sky130_fd_sc_hd__inv_1
X$8064 \$153 \$9406 \$9252 \$9324 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8065 \$153 \$9407 \$8917 \$9276 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8067 \$16 \$8220 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8068 \$16 \$7709 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8070 \$153 \$9360 \$9278 \$8891 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8071 \$16 \$8220 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8072 \$16 \$9253 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8073 \$153 \$9429 \$9081 \$9253 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8074 \$153 \$9277 \$9081 \$9214 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8075 \$16 \$8044 \$9518 \$9431 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$8078 \$153 \$9430 \$9133 \$9276 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8079 \$16 \$9214 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8080 \$153 \$9375 \$8937 \$9253 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8082 \$153 \$9375 \$9252 \$8843 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8083 \$153 \$9250 \$8917 \$7994 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8085 \$153 \$9303 \$8917 \$8993 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8087 \$16 \$8936 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8088 \$153 \$9432 \$9174 \$9325 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8089 \$153 \$9345 \$9466 \$8936 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8090 \$153 \$9466 \$8772 \$9305 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$8091 \$153 \$9433 \$7915 \$9520 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$8094 \$153 \$9387 \$8842 \$9521 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8095 \$153 \$9306 \$9047 \$9033 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8096 \$16 \$7691 \$16 \$153 \$9521 VNB sky130_fd_sc_hd__inv_1
X$8097 \$16 \$7691 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8098 \$16 \$8807 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8099 \$153 \$9434 \$9408 \$8807 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8101 \$153 \$9435 \$8842 \$9409 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8103 \$16 \$7695 \$16 \$153 \$9409 VNB sky130_fd_sc_hd__inv_1
X$8105 \$16 \$7695 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8106 \$153 \$9408 \$8101 \$9436 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$8107 \$16 \$7695 \$8960 \$9436 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$8108 \$153 \$9437 \$9347 \$9253 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8109 \$153 \$9231 \$8917 \$9151 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8110 \$153 \$9437 \$9252 \$9328 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8113 \$153 \$9376 \$9347 \$9275 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8114 \$153 \$9376 \$9278 \$9328 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8115 \$153 \$9467 \$7852 \$9438 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$8116 \$16 \$7347 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8118 \$16 \$7793 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8119 \$16 \$7793 \$16 \$153 \$9439 VNB sky130_fd_sc_hd__inv_1
X$8120 \$153 \$9410 \$9256 \$9439 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8122 \$153 \$9440 \$8996 \$9439 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8124 \$16 \$9035 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8125 \$16 \$7344 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8127 \$153 \$9263 \$9179 \$9034 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8128 \$16 \$9034 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8129 \$16 \$7709 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8130 \$16 \$7903 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8131 \$153 \$9441 \$7903 \$9388 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$8132 \$16 \$7709 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8133 \$16 \$7709 \$16 \$153 \$9329 VNB sky130_fd_sc_hd__inv_1
X$8135 \$153 \$9351 \$9441 \$9034 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8136 \$153 \$9456 \$9441 \$8927 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8137 \$153 \$9377 \$9279 \$9134 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8138 \$16 \$8893 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8139 \$16 \$9191 \$16 \$153 \$9675 VNB sky130_fd_sc_hd__clkbuf_2
X$8140 \$16 \$9034 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8142 \$153 \$9378 \$9279 \$9034 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8143 \$153 \$9378 \$9059 \$9264 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8144 \$153 \$9379 \$9279 \$8844 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8145 \$153 \$9379 \$8965 \$9264 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8146 \$16 \$7691 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8147 \$16 \$9191 \$16 \$153 \$8825 VNB sky130_fd_sc_hd__clkbuf_2
X$8149 \$153 \$9389 \$8977 \$9411 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8151 \$16 \$7915 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8152 \$16 \$7691 \$8825 \$9442 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$8153 \$153 \$9364 \$7915 \$9442 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$8155 \$153 \$9281 \$9364 \$9134 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8156 \$16 \$9134 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8158 \$16 \$7691 \$16 \$153 \$9280 VNB sky130_fd_sc_hd__inv_1
X$8159 \$16 \$8893 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8161 \$153 \$9443 \$9364 \$8893 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8162 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$8163 \$16 \$8927 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8164 \$153 \$9380 \$9316 \$8927 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8165 \$153 \$9444 \$9316 \$9034 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8166 \$16 \$9034 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8169 \$16 \$7695 \$8825 \$9390 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$8170 \$153 \$9391 \$8101 \$9390 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$8171 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$8172 \$16 \$9134 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8173 \$153 \$9446 \$9391 \$9134 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8174 \$153 \$9445 \$8996 \$9366 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8176 \$16 \$9034 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8178 \$153 \$9282 \$9240 \$9034 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8179 \$153 \$9447 \$9391 \$9154 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8181 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$8182 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$8183 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$8185 \$153 \$1091 \$1036 \$17 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8187 \$153 \$1091 \$102 \$1012 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8188 \$153 \$1137 \$561 \$1012 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8190 \$16 \$783 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8191 \$153 \$1116 \$30 \$1012 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8194 \$153 \$1092 \$1036 \$249 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8195 \$153 \$1092 \$377 \$1012 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8196 \$153 \$951 \$1036 \$419 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8197 \$153 \$1065 \$59 \$1012 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8198 \$16 \$184 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8199 \$16 \$419 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8200 \$16 \$981 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8202 \$153 \$1125 \$59 \$1106 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8203 \$153 \$1429 \$561 \$1106 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8204 \$153 \$663 \$952 \$504 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8205 \$16 \$504 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8206 \$16 \$537 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8207 \$153 \$1066 \$394 \$903 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8208 \$153 \$1107 \$561 \$903 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8211 \$153 \$922 \$377 \$903 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8212 \$153 \$923 \$349 \$903 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8213 \$153 \$1093 \$817 \$263 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8214 \$153 \$1019 \$59 \$639 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8215 \$153 \$1093 \$234 \$639 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8216 \$16 \$1067 \$16 \$153 \$639 VNB sky130_fd_sc_hd__inv_1
X$8218 \$153 \$1117 \$394 \$1191 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8219 \$16 \$537 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8221 \$153 \$1126 \$1118 \$17 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8222 \$16 \$263 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8224 \$153 \$1138 \$1118 \$184 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8225 \$153 \$1108 \$30 \$1193 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8227 \$16 \$184 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8228 \$16 \$249 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8230 \$153 \$1108 \$1118 \$58 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8231 \$153 \$975 \$394 \$651 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8232 \$16 \$58 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8234 \$153 \$1127 \$1038 \$263 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8235 \$16 \$395 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8236 \$16 \$263 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8237 \$16 \$17 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8240 \$153 \$1094 \$1038 \$58 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8241 \$153 \$1094 \$30 \$1070 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8242 \$153 \$1095 \$955 \$419 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8243 \$153 \$1095 \$349 \$906 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8244 \$16 \$249 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8245 \$16 \$58 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8246 \$16 \$58 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8248 \$16 \$184 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8249 \$16 \$715 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8251 \$16 \$1048 \$16 \$153 \$906 VNB sky130_fd_sc_hd__inv_1
X$8252 \$153 \$978 \$102 \$906 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8253 \$153 \$1071 \$394 \$906 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8254 \$16 \$1037 \$979 \$1072 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$8255 \$153 \$1096 \$1039 \$209 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8256 \$153 \$1096 \$346 \$1196 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8258 \$153 \$1128 \$1039 \$73 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8259 \$16 \$73 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8261 \$153 \$1174 \$1039 \$60 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8262 \$153 \$1097 \$1039 \$18 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8264 \$16 \$981 \$16 \$153 \$767 VNB sky130_fd_sc_hd__inv_1
X$8266 \$153 \$1075 \$347 \$767 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8267 \$16 \$1013 \$507 \$1175 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$8268 \$16 \$507 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8269 \$153 \$1129 \$956 \$209 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8270 \$153 \$1109 \$35 \$767 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8271 \$16 \$60 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8272 \$16 \$212 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8273 \$16 \$1067 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8276 \$16 \$1211 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8277 \$153 \$1076 \$215 \$1111 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8278 \$16 \$209 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8279 \$153 \$1110 \$823 \$209 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8280 \$153 \$1049 \$347 \$1111 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8281 \$153 \$983 \$54 \$1111 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8282 \$16 \$1067 \$507 \$1130 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$8283 \$16 \$293 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8286 \$16 \$908 \$16 \$153 \$507 VNB sky130_fd_sc_hd__clkbuf_2
X$8287 \$153 \$1098 \$900 \$293 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8288 \$153 \$1098 \$35 \$909 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8289 \$16 \$1067 \$16 \$153 \$909 VNB sky130_fd_sc_hd__inv_1
X$8291 \$153 \$988 \$253 \$909 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8292 \$153 \$1110 \$346 \$1040 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8293 \$16 \$358 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8295 \$16 \$293 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8297 \$153 \$1112 \$1041 \$187 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8298 \$153 \$1077 \$104 \$1199 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8299 \$16 \$187 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8300 \$153 \$1140 \$957 \$187 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8301 \$153 \$1112 \$54 \$1199 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8302 \$16 \$187 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8303 \$16 \$358 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8305 \$153 \$1141 \$957 \$209 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8306 \$16 \$1551 \$946 \$1131 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$8308 \$153 \$1142 \$1042 \$60 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8309 \$153 \$1050 \$1042 \$187 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8310 \$16 \$209 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8312 \$153 \$1143 \$1042 \$212 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8313 \$153 \$1080 \$346 \$1051 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8314 \$153 \$1132 \$1026 \$241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8315 \$153 \$993 \$21 \$947 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8316 \$16 \$424 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8318 \$16 \$79 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8320 \$153 \$1052 \$1026 \$79 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8322 \$16 \$1489 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8323 \$153 \$1082 \$44 \$947 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8325 \$16 \$902 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8326 \$153 \$994 \$353 \$657 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8328 \$16 \$82 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8330 \$16 \$2232 \$268 \$1113 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$8331 \$153 \$854 \$1245 \$1113 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$8332 \$153 \$1144 \$958 \$424 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8334 \$16 \$798 \$16 \$153 \$813 VNB sky130_fd_sc_hd__inv_1
X$8335 \$153 \$958 \$856 \$1054 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$8336 \$153 \$1145 \$958 \$145 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8337 \$16 \$1201 \$16 \$153 \$268 VNB sky130_fd_sc_hd__clkbuf_2
X$8338 \$16 \$145 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8342 \$16 \$82 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8344 \$16 \$424 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8345 \$16 \$79 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8346 \$153 \$1135 \$1056 \$79 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8347 \$153 \$1146 \$1056 \$424 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8348 \$153 \$1084 \$389 \$814 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8349 \$16 \$273 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8350 \$16 \$2462 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8353 \$16 \$1719 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8354 \$16 \$79 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8355 \$16 \$145 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8356 \$153 \$1101 \$1043 \$79 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8357 \$153 \$1101 \$112 \$1057 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8358 \$153 \$1114 \$559 \$1456 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8360 \$153 \$1102 \$893 \$82 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8361 \$153 \$1375 \$353 \$1205 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8362 \$153 \$1102 \$44 \$915 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8364 \$153 \$893 \$1303 \$1119 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$8365 \$16 \$1120 \$441 \$1119 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$8366 \$16 \$1121 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8368 \$16 \$441 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8369 \$16 \$1120 \$16 \$153 \$915 VNB sky130_fd_sc_hd__inv_1
X$8370 \$153 \$1086 \$388 \$915 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8371 \$153 \$1319 \$559 \$1811 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8372 \$16 \$446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8373 \$16 \$178 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8374 \$153 \$1103 \$1058 \$178 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8375 \$153 \$1103 \$549 \$1087 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8376 \$16 \$149 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8377 \$16 \$509 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8379 \$153 \$1122 \$393 \$1087 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8381 \$153 \$1104 \$1058 \$509 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8382 \$153 \$1104 \$371 \$1087 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8383 \$153 \$1147 \$1245 \$1123 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$8385 \$16 \$423 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8387 \$153 \$1148 \$1147 \$309 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8388 \$153 \$1124 \$371 \$1059 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8389 \$16 \$1062 \$16 \$153 \$615 VNB sky130_fd_sc_hd__clkbuf_2
X$8390 \$153 \$942 \$57 \$659 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8391 \$16 \$615 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8393 \$16 \$1062 \$16 \$153 \$428 VNB sky130_fd_sc_hd__clkbuf_2
X$8394 \$16 \$2462 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8395 \$16 \$178 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8396 \$153 \$1105 \$1278 \$178 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8397 \$153 \$1105 \$549 \$1115 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8399 \$153 \$1149 \$1006 \$446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8400 \$16 \$1184 \$16 \$153 \$949 VNB sky130_fd_sc_hd__inv_1
X$8402 \$16 \$178 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8404 \$153 \$1150 \$1006 \$178 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8405 \$153 \$1151 \$1006 \$63 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8406 \$153 \$1280 \$1006 \$509 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8407 \$16 \$509 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8409 \$16 \$815 \$16 \$153 \$776 VNB sky130_fd_sc_hd__inv_1
X$8410 \$16 \$309 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8412 \$153 \$1152 \$943 \$309 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8413 \$153 \$1088 \$549 \$776 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8414 \$16 \$63 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8415 \$153 \$1136 \$966 \$309 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8416 \$153 \$1089 \$57 \$898 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8417 \$16 \$309 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8418 \$16 \$1228 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8420 \$16 \$1120 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8421 \$16 \$895 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8423 \$16 \$446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8424 \$16 \$310 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8425 \$153 \$1010 \$549 \$898 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8427 \$153 \$1153 \$1186 \$310 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8428 \$153 \$1090 \$393 \$898 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8429 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$8431 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$8432 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$8433 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$8434 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$8435 \$153 \$1137 \$1036 \$504 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8436 \$16 \$504 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8437 \$16 \$17 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8440 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$8441 \$153 \$1116 \$1036 \$58 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8442 \$16 \$58 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8443 \$16 \$58 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8444 \$16 \$783 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8445 \$16 \$1168 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8446 \$153 \$1207 \$377 \$1187 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8448 \$16 \$1037 \$1168 \$1064 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$8449 \$153 \$1036 \$1208 \$1169 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$8451 \$16 \$981 \$1168 \$1169 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$8452 \$153 \$1125 \$1257 \$184 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8454 \$153 \$1188 \$30 \$1106 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8455 \$153 \$1154 \$952 \$58 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8456 \$153 \$1154 \$30 \$783 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8458 \$16 \$1291 \$16 \$153 \$783 VNB sky130_fd_sc_hd__inv_1
X$8459 \$153 \$1189 \$102 \$783 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8460 \$16 \$1013 \$537 \$1209 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$8462 \$153 \$1107 \$755 \$504 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8463 \$16 \$1013 \$16 \$153 \$903 VNB sky130_fd_sc_hd__inv_1
X$8464 \$16 \$504 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8466 \$16 \$537 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8467 \$153 \$817 \$1211 \$1170 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$8469 \$16 \$1067 \$537 \$1170 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$8471 \$16 \$263 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8472 \$153 \$1117 \$1258 \$395 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8474 \$153 \$1190 \$561 \$1191 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8475 \$16 \$1192 \$16 \$153 \$1168 VNB sky130_fd_sc_hd__clkbuf_2
X$8476 \$16 \$395 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8477 \$153 \$1210 \$1118 \$263 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8479 \$153 \$1126 \$102 \$1193 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8480 \$16 \$1211 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8481 \$153 \$1212 \$1118 \$249 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8482 \$16 \$691 \$715 \$1213 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$8484 \$153 \$1172 \$1118 \$395 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8485 \$16 \$395 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8486 \$16 \$715 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8487 \$16 \$1171 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8491 \$16 \$715 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8492 \$153 \$1155 \$1038 \$395 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8493 \$153 \$1022 \$561 \$1193 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8494 \$153 \$1172 \$394 \$1193 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8495 \$153 \$1194 \$59 \$1070 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8496 \$153 \$977 \$377 \$1070 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8499 \$153 \$1214 \$955 \$249 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8500 \$16 \$1182 \$1332 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$8501 \$16 \$1407 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8502 \$153 \$1156 \$955 \$58 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8503 \$153 \$1156 \$30 \$906 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8504 \$153 \$1195 \$59 \$906 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8507 \$153 \$1157 \$1039 \$187 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8508 \$153 \$1157 \$54 \$1196 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8509 \$16 \$1390 \$16 \$153 \$1196 VNB sky130_fd_sc_hd__inv_1
X$8510 \$16 \$209 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8512 \$153 \$1128 \$215 \$1196 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8513 \$153 \$1215 \$1039 \$212 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8516 \$153 \$1174 \$104 \$1196 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8517 \$153 \$758 \$1208 \$1216 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$8518 \$153 \$1109 \$758 \$293 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8520 \$153 \$956 \$972 \$1175 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$8523 \$153 \$1217 \$956 \$60 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8525 \$153 \$1218 \$956 \$18 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8526 \$16 \$1291 \$507 \$1197 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$8527 \$16 \$18 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8528 \$153 \$1158 \$823 \$212 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8530 \$153 \$1159 \$823 \$293 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8531 \$153 \$900 \$1211 \$1130 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$8532 \$153 \$1160 \$900 \$187 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8533 \$153 \$1160 \$54 \$909 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8536 \$16 \$187 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8537 \$153 \$1198 \$347 \$909 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8538 \$153 \$1219 \$1041 \$293 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8540 \$153 \$1220 \$1041 \$212 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8541 \$153 \$1078 \$215 \$1199 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8542 \$16 \$212 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8545 \$153 \$1221 \$957 \$293 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8546 \$16 \$1048 \$16 \$153 \$910 VNB sky130_fd_sc_hd__inv_1
X$8548 \$153 \$1176 \$957 \$212 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8549 \$153 \$1141 \$346 \$910 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8550 \$153 \$1176 \$347 \$910 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8551 \$16 \$293 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8553 \$153 \$1177 \$35 \$1051 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8554 \$153 \$1142 \$104 \$1051 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8555 \$153 \$1200 \$215 \$1411 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8556 \$153 \$1222 \$1042 \$358 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8558 \$153 \$1143 \$347 \$1051 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8560 \$16 \$21 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8562 \$153 \$1161 \$1026 \$424 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8563 \$153 \$1161 \$353 \$947 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8565 \$153 \$1081 \$266 \$947 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8567 \$153 \$1026 \$1489 \$1223 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$8568 \$16 \$1044 \$16 \$153 \$947 VNB sky130_fd_sc_hd__inv_1
X$8571 \$16 \$79 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8572 \$153 \$1224 \$1183 \$79 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8573 \$16 \$1044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8575 \$16 \$2232 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8576 \$16 \$79 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8577 \$153 \$1225 \$854 \$79 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8578 \$153 \$1083 \$44 \$657 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8579 \$16 \$2232 \$16 \$153 \$657 VNB sky130_fd_sc_hd__inv_1
X$8582 \$153 \$1134 \$21 \$657 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8584 \$153 \$1053 \$958 \$241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8585 \$153 \$1144 \$353 \$813 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8587 \$16 \$1201 \$16 \$153 \$397 VNB sky130_fd_sc_hd__clkbuf_2
X$8588 \$153 \$1055 \$958 \$79 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8591 \$153 \$1145 \$266 \$813 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8592 \$16 \$1201 \$16 \$153 \$441 VNB sky130_fd_sc_hd__clkbuf_2
X$8594 \$153 \$1202 \$1056 \$241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8595 \$153 \$1162 \$1056 \$82 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8596 \$153 \$1202 \$388 \$814 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8598 \$153 \$1162 \$44 \$814 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8599 \$153 \$1146 \$353 \$814 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8600 \$16 \$2462 \$16 \$153 \$814 VNB sky130_fd_sc_hd__inv_1
X$8601 \$153 \$1163 \$1043 \$273 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8602 \$153 \$1163 \$389 \$1057 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8603 \$153 \$1203 \$353 \$1057 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8606 \$16 \$1184 \$16 \$153 \$1057 VNB sky130_fd_sc_hd__inv_1
X$8608 \$16 \$82 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8609 \$153 \$1227 \$1185 \$82 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8610 \$16 \$82 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8612 \$153 \$1204 \$389 \$1205 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8613 \$16 \$79 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8614 \$16 \$273 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8615 \$16 \$1228 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8617 \$153 \$882 \$559 \$915 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8618 \$153 \$1085 \$112 \$915 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8619 \$153 \$1398 \$112 \$1229 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8621 \$16 \$1044 \$369 \$1230 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$8622 \$153 \$1178 \$266 \$1205 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8623 \$153 \$1058 \$1489 \$1230 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$8625 \$153 \$1122 \$1058 \$446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8626 \$153 \$1231 \$1058 \$63 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8627 \$16 \$63 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8629 \$16 \$309 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8630 \$16 \$310 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8631 \$153 \$1164 \$1058 \$310 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8634 \$153 \$1164 \$223 \$1087 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8635 \$16 \$2232 \$428 \$1123 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$8636 \$16 \$964 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8637 \$16 \$149 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8638 \$153 \$1060 \$1147 \$149 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8639 \$16 \$2232 \$16 \$153 \$1059 VNB sky130_fd_sc_hd__inv_1
X$8640 \$16 \$309 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8641 \$153 \$1124 \$1147 \$509 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8644 \$153 \$1148 \$703 \$1059 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8645 \$16 \$2462 \$615 \$1232 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$8646 \$153 \$1063 \$1278 \$310 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8647 \$16 \$310 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8649 \$16 \$509 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8650 \$16 \$309 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8651 \$153 \$1233 \$1278 \$309 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8653 \$16 \$1719 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8656 \$153 \$1006 \$1719 \$1179 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$8657 \$16 \$1184 \$615 \$1179 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$8659 \$153 \$1149 \$393 \$949 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8660 \$16 \$309 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8661 \$153 \$1150 \$549 \$949 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8663 \$16 \$63 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8665 \$16 \$310 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8667 \$153 \$1151 \$57 \$949 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8669 \$153 \$1165 \$943 \$310 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8670 \$153 \$1165 \$223 \$776 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8672 \$16 \$1120 \$615 \$1181 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$8673 \$153 \$966 \$1303 \$1181 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$8676 \$153 \$1166 \$1186 \$509 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8677 \$153 \$1166 \$371 \$1206 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8678 \$16 \$149 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8679 \$153 \$1167 \$1186 \$149 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8680 \$153 \$1167 \$398 \$1206 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8681 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$8683 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$8685 \$153 \$1153 \$223 \$1206 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8686 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$8687 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$8688 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$8689 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$8690 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$8692 \$153 \$1282 \$1256 \$504 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8693 \$16 \$504 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8694 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$8696 \$153 \$1234 \$1256 \$58 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8697 \$153 \$1234 \$30 \$1187 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8701 \$16 \$1037 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8702 \$153 \$1235 \$1256 \$419 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8703 \$153 \$1235 \$349 \$1187 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8704 \$16 \$419 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8706 \$16 \$1168 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8707 \$153 \$1188 \$1257 \$58 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8708 \$16 \$58 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8709 \$16 \$1208 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8710 \$16 \$981 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8714 \$16 \$754 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8715 \$153 \$1046 \$952 \$249 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8716 \$153 \$1189 \$952 \$17 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8718 \$153 \$755 \$972 \$1209 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$8719 \$16 \$1291 \$537 \$1283 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$8722 \$16 \$1522 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8723 \$16 \$537 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8724 \$16 \$541 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8726 \$153 \$1236 \$1249 \$17 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8727 \$153 \$1236 \$102 \$1250 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8728 \$16 \$17 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8729 \$16 \$17 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8730 \$153 \$1237 \$1258 \$17 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8731 \$16 \$1192 \$16 \$153 \$537 VNB sky130_fd_sc_hd__clkbuf_2
X$8733 \$153 \$1237 \$102 \$1191 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8734 \$16 \$1192 \$16 \$153 \$503 VNB sky130_fd_sc_hd__clkbuf_2
X$8736 \$153 \$1284 \$1118 \$419 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8737 \$16 \$419 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8738 \$16 \$395 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8739 \$16 \$1067 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8740 \$153 \$1212 \$377 \$1193 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8741 \$153 \$1138 \$59 \$1193 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8742 \$16 \$263 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8744 \$153 \$1118 \$842 \$1213 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$8745 \$16 \$691 \$16 \$153 \$1193 VNB sky130_fd_sc_hd__inv_1
X$8746 \$16 \$715 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8747 \$16 \$715 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8749 \$153 \$1259 \$234 \$1251 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8751 \$153 \$1285 \$1038 \$17 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8752 \$16 \$184 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8753 \$16 \$1331 \$505 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$8754 \$16 \$1331 \$541 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$8756 \$153 \$1194 \$1038 \$184 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8757 \$16 \$1331 \$972 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$8758 \$16 \$1048 \$715 \$1260 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$8759 \$153 \$955 \$1173 \$1260 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$8760 \$16 \$1182 \$1173 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$8761 \$153 \$1214 \$377 \$906 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8762 \$16 \$1182 \$1139 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$8763 \$16 \$16 \$153 VNB sky130_fd_sc_hd__conb_1
X$8765 \$153 \$1195 \$955 \$184 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8766 \$153 \$382 \$394 \$173 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8768 \$153 \$1287 \$1261 \$293 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8769 \$16 \$293 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8770 \$153 \$1073 \$35 \$1196 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8771 \$16 \$187 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8774 \$153 \$1287 \$35 \$1409 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8776 \$16 \$73 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8777 \$153 \$1074 \$253 \$1196 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8779 \$153 \$1288 \$1261 \$18 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8780 \$153 \$1215 \$347 \$1196 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8781 \$16 \$981 \$979 \$1216 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$8782 \$16 \$18 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8785 \$153 \$1289 \$1262 \$293 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8786 \$16 \$293 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8788 \$153 \$1290 \$1262 \$18 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8789 \$16 \$18 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8790 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$8791 \$16 \$1291 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8792 \$153 \$1217 \$104 \$1111 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8793 \$16 \$1013 \$16 \$153 \$1111 VNB sky130_fd_sc_hd__inv_1
X$8794 \$16 \$1013 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8796 \$16 \$1263 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8797 \$16 \$507 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8798 \$153 \$823 \$1263 \$1197 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$8800 \$16 \$1292 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8801 \$16 \$212 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8802 \$16 \$1291 \$16 \$153 \$1040 VNB sky130_fd_sc_hd__inv_1
X$8803 \$153 \$1265 \$823 \$187 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8804 \$16 \$908 \$16 \$153 \$979 VNB sky130_fd_sc_hd__clkbuf_2
X$8807 \$153 \$985 \$104 \$1040 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8808 \$153 \$1198 \$900 \$212 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8809 \$16 \$212 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8811 \$153 \$1293 \$1041 \$18 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8812 \$16 \$1264 \$16 \$153 \$1199 VNB sky130_fd_sc_hd__inv_1
X$8814 \$153 \$1265 \$54 \$1040 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8816 \$16 \$1048 \$946 \$1266 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$8817 \$153 \$957 \$1173 \$1266 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$8818 \$153 \$1220 \$347 \$1199 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8819 \$153 \$1219 \$35 \$1199 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8820 \$153 \$1140 \$54 \$910 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8822 \$16 \$293 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8823 \$153 \$1042 \$1139 \$1131 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$8824 \$16 \$212 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8825 \$153 \$1177 \$1042 \$293 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8826 \$153 \$1295 \$1336 \$209 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8827 \$16 \$1551 \$16 \$153 \$1051 VNB sky130_fd_sc_hd__inv_1
X$8829 \$16 \$73 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8831 \$153 \$1317 \$1042 \$73 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8832 \$16 \$358 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8833 \$16 \$1551 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8834 \$16 \$273 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8835 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8836 \$153 \$1294 \$1482 \$21 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8837 \$153 \$1296 \$1026 \$273 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8839 \$153 \$153 \$353 \$1337 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8840 \$16 \$1044 \$397 \$1223 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$8842 \$16 \$82 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8843 \$153 \$1297 \$1183 \$82 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8844 \$16 \$397 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8845 \$16 \$1044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8847 \$16 \$2232 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8849 \$153 \$1133 \$559 \$657 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8850 \$16 \$265 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8851 \$153 \$1298 \$1268 \$79 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8852 \$153 \$1224 \$112 \$1252 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8854 \$153 \$1269 \$21 \$1396 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8855 \$16 \$1433 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8856 \$16 \$1433 \$16 \$153 \$1201 VNB sky130_fd_sc_hd__clkbuf_2
X$8857 \$153 \$741 \$559 \$913 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8858 \$153 \$857 \$44 \$913 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8859 \$16 \$241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8860 \$16 \$79 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8862 \$16 \$79 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8865 \$153 \$1239 \$1270 \$79 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8866 \$16 \$268 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8867 \$153 \$1056 \$1272 \$1271 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$8868 \$153 \$1300 \$1254 \$79 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8869 \$16 \$79 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8870 \$16 \$1272 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8872 \$16 \$424 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8874 \$153 \$1203 \$1043 \$424 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8875 \$153 \$1043 \$1719 \$1273 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$8876 \$16 \$1184 \$441 \$1273 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$8877 \$153 \$1226 \$559 \$1057 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8878 \$153 \$1274 \$21 \$1240 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8881 \$153 \$1204 \$1185 \$273 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8883 \$16 \$1228 \$441 \$1241 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$8884 \$153 \$1301 \$1185 \$79 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8885 \$153 \$1185 \$1121 \$1241 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$8886 \$16 \$145 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8887 \$16 \$241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8889 \$153 \$1242 \$1185 \$241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8890 \$153 \$1242 \$388 \$1205 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8891 \$16 \$1228 \$16 \$153 \$1205 VNB sky130_fd_sc_hd__inv_1
X$8893 \$153 \$153 \$549 \$1243 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8894 \$153 \$153 \$703 \$1243 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8895 \$153 \$153 \$371 \$1243 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8897 \$153 \$1231 \$57 \$1087 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8898 \$153 \$1244 \$1058 \$309 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8899 \$153 \$1244 \$703 \$1087 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8901 \$16 \$1245 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8902 \$153 \$1275 \$549 \$1341 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8903 \$16 \$310 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8904 \$16 \$428 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8905 \$16 \$265 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8906 \$16 \$2232 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8907 \$16 \$399 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8909 \$16 \$2232 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8910 \$16 \$509 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8911 \$153 \$1276 \$223 \$1059 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8912 \$153 \$1277 \$549 \$1059 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8913 \$16 \$1272 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8914 \$16 \$149 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8915 \$153 \$1278 \$1272 \$1232 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$8916 \$153 \$1246 \$1278 \$149 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8918 \$153 \$1246 \$398 \$1115 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8919 \$153 \$1247 \$1278 \$509 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8920 \$153 \$1233 \$703 \$1115 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8921 \$153 \$1247 \$371 \$1115 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8922 \$16 \$615 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8923 \$16 \$1184 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8924 \$153 \$1279 \$398 \$1255 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8926 \$16 \$1184 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8927 \$16 \$149 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8929 \$153 \$1248 \$1302 \$149 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8930 \$153 \$1280 \$371 \$949 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8931 \$153 \$1248 \$398 \$1343 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8932 \$16 \$1120 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8933 \$16 \$1303 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8934 \$16 \$615 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8935 \$16 \$1121 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8937 \$16 \$509 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8938 \$153 \$1152 \$703 \$776 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8939 \$153 \$1186 \$1121 \$1281 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$8940 \$153 \$1304 \$1186 \$63 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8941 \$16 \$509 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8942 \$153 \$1304 \$57 \$1206 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8943 \$16 \$1228 \$16 \$153 \$1206 VNB sky130_fd_sc_hd__inv_1
X$8946 \$153 \$1305 \$1186 \$178 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8948 \$153 \$1307 \$1186 \$446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8949 \$16 \$446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8950 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$8952 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$8953 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$8954 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$8955 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$8957 \$153 \$1045 \$1036 \$263 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8958 \$16 \$263 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8959 \$16 \$17 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8962 \$153 \$1282 \$561 \$1187 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8963 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$8964 \$153 \$1207 \$1256 \$249 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8965 \$16 \$249 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8966 \$16 \$1390 \$1168 \$1310 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$8967 \$153 \$1256 \$1311 \$1310 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$8968 \$16 \$1390 \$16 \$153 \$1187 VNB sky130_fd_sc_hd__inv_1
X$8969 \$16 \$1168 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8970 \$16 \$1037 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8972 \$16 \$1311 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8973 \$16 \$1390 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8974 \$153 \$1312 \$1257 \$17 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8975 \$16 \$17 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8976 \$153 \$1312 \$102 \$1106 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8977 \$153 \$1313 \$1326 \$504 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8978 \$153 \$1313 \$561 \$1327 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8980 \$16 \$17 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8982 \$16 \$17 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8983 \$153 \$952 \$1263 \$1283 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$8984 \$153 \$1346 \$1249 \$419 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8986 \$153 \$1347 \$1249 \$263 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8987 \$16 \$419 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8988 \$16 \$263 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8990 \$16 \$1328 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8991 \$16 \$1328 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8992 \$16 \$1168 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8993 \$16 \$1348 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8994 \$153 \$1190 \$1258 \$504 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$8996 \$153 \$1329 \$349 \$1191 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$8997 \$16 \$504 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$8998 \$16 \$1192 \$16 \$153 \$715 VNB sky130_fd_sc_hd__clkbuf_2
X$8999 \$153 \$1452 \$1330 \$395 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9001 \$153 \$1349 \$1330 \$263 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9002 \$16 \$1551 \$715 \$1350 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$9003 \$153 \$1352 \$1171 \$1351 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$9004 \$153 \$1259 \$1352 \$263 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9005 \$16 \$263 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9006 \$16 \$17 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9009 \$153 \$1353 \$1352 \$504 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9010 \$153 \$1389 \$394 \$1251 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9011 \$153 \$1285 \$102 \$1070 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9012 \$16 \$1331 \$684 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$9013 \$16 \$1508 \$715 \$1314 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$9014 \$153 \$1038 \$1332 \$1314 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$9016 \$153 \$1069 \$561 \$1070 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9017 \$16 \$1182 \$685 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$9018 \$16 \$1182 \$1171 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$9019 \$16 \$1182 \$584 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$9020 \$16 \$1182 \$842 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$9021 \$153 \$153 \$561 \$1408 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9022 \$153 \$153 \$234 \$1408 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9023 \$16 \$1354 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9024 \$153 \$1039 \$1311 \$1355 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$9027 \$153 \$1308 \$1261 \$209 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9028 \$16 \$209 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9029 \$16 \$187 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9030 \$16 \$1311 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9031 \$153 \$1356 \$1261 \$73 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9032 \$153 \$1469 \$1261 \$358 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9033 \$16 \$358 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9035 \$153 \$1357 \$1261 \$60 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9036 \$16 \$60 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9037 \$16 \$18 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9039 \$16 \$979 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9040 \$153 \$1315 \$1262 \$187 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9041 \$153 \$1315 \$54 \$1333 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9042 \$16 \$187 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9043 \$16 \$358 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9044 \$16 \$293 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9048 \$153 \$1391 \$253 \$1333 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9049 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$9051 \$153 \$1358 \$1334 \$73 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9052 \$153 \$1129 \$346 \$1111 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9053 \$153 \$984 \$35 \$1111 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9054 \$16 \$73 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9055 \$16 \$358 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9057 \$153 \$1359 \$253 \$1393 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9058 \$16 \$187 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9059 \$153 \$1316 \$1421 \$18 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9060 \$153 \$1014 \$215 \$1040 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9061 \$16 \$18 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9062 \$153 \$1360 \$215 \$1335 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9064 \$16 \$1067 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9066 \$16 \$1264 \$946 \$1395 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$9067 \$153 \$1361 \$1041 \$358 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9068 \$153 \$1362 \$1041 \$209 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9069 \$16 \$209 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9070 \$153 \$1336 \$1332 \$1363 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$9072 \$153 \$1364 \$1336 \$358 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9073 \$153 \$1221 \$35 \$910 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9074 \$153 \$1364 \$253 \$1411 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9075 \$16 \$358 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9076 \$153 \$1365 \$1336 \$293 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9077 \$16 \$293 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9078 \$16 \$60 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9080 \$153 \$1366 \$1336 \$60 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9082 \$153 \$1516 \$18 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$9083 \$16 \$1516 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9085 \$153 \$1317 \$215 \$1051 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9086 \$16 \$1406 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9087 \$16 \$1811 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9088 \$16 \$1367 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9092 \$16 \$1538 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9093 \$153 \$1538 \$79 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$9094 \$153 \$1296 \$389 \$947 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9095 \$16 \$16 \$153 VNB sky130_fd_sc_hd__conb_1
X$9096 \$16 \$1378 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9097 \$153 \$153 \$559 \$1337 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9098 \$153 \$153 \$389 \$1337 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9101 \$16 \$273 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9103 \$153 \$1027 \$266 \$657 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9104 \$16 \$1245 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9105 \$16 \$268 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9106 \$16 \$964 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9107 \$16 \$79 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9109 \$153 \$1297 \$44 \$1252 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9110 \$16 \$241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9111 \$16 \$79 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9113 \$16 \$82 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9114 \$16 \$79 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9116 \$153 \$1370 \$1253 \$79 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9118 \$16 \$2462 \$441 \$1271 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$9120 \$153 \$1135 \$112 \$814 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9121 \$153 \$1339 \$44 \$1412 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9122 \$16 \$441 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9123 \$16 \$79 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9124 \$153 \$1372 \$1320 \$79 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9127 \$153 \$1373 \$266 \$1240 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9128 \$153 \$1374 \$559 \$1240 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9130 \$16 \$273 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9131 \$153 \$1375 \$1185 \$424 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9133 \$153 \$1227 \$44 \$1205 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9134 \$153 \$1301 \$112 \$1205 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9135 \$153 \$1178 \$1185 \$145 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9136 \$16 \$1378 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9137 \$16 \$369 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9139 \$16 \$16 \$153 VNB sky130_fd_sc_hd__conb_1
X$9140 \$16 \$1228 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9141 \$153 \$153 \$23 \$1243 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9142 \$153 \$153 \$393 \$1243 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9144 \$16 \$309 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9145 \$153 \$1322 \$1340 \$309 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9146 \$153 \$1322 \$703 \$1341 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9147 \$16 \$964 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9149 \$16 \$178 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9151 \$153 \$1275 \$1340 \$178 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9153 \$153 \$1276 \$1147 \$310 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9154 \$16 \$178 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9155 \$16 \$258 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9157 \$16 \$446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9158 \$153 \$1323 \$1147 \$446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9160 \$153 \$1323 \$393 \$1059 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9161 \$16 \$1485 \$16 \$153 \$1062 VNB sky130_fd_sc_hd__clkbuf_2
X$9162 \$153 \$1380 \$1278 \$446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9163 \$153 \$1379 \$23 \$1115 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9164 \$16 \$901 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9166 \$16 \$2462 \$16 \$153 \$1115 VNB sky130_fd_sc_hd__inv_1
X$9167 \$16 \$2462 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9168 \$153 \$1478 \$1342 \$310 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9170 \$153 \$1382 \$1302 \$310 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9173 \$153 \$1383 \$23 \$1343 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9174 \$16 \$815 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9175 \$16 \$63 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9176 \$153 \$1384 \$943 \$63 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9177 \$153 \$1385 \$943 \$509 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9178 \$16 \$1228 \$615 \$1281 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$9179 \$16 \$63 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9181 \$16 \$309 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9183 \$153 \$1324 \$1186 \$309 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9184 \$153 \$1324 \$703 \$1206 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9185 \$153 \$1386 \$57 \$1344 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9186 \$16 \$178 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9187 \$153 \$1305 \$549 \$1206 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9188 \$153 \$1387 \$703 \$1344 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9191 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$9193 \$153 \$1306 \$23 \$1206 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9194 \$153 \$1345 \$223 \$1415 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9195 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$9196 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$9197 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$9199 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$9200 \$153 \$8360 \$8331 \$6981 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9201 \$153 \$8431 \$6749 \$8384 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9202 \$16 \$6981 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9204 \$153 \$8406 \$8331 \$6907 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9205 \$153 \$8406 \$6913 \$8384 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9207 \$16 \$8139 \$8024 \$8456 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$9208 \$153 \$8432 \$6719 \$8384 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9209 \$16 \$6792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9211 \$153 \$8433 \$8333 \$6860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9212 \$153 \$8433 \$6732 \$8206 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9213 \$153 \$8434 \$8638 \$7816 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9214 \$16 \$8423 \$8024 \$8421 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$9216 \$153 \$8435 \$8912 \$7816 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9217 \$153 \$8407 \$8115 \$7041 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9218 \$153 \$8407 \$6996 \$8036 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9219 \$16 \$7041 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9220 \$16 \$8271 \$8024 \$8408 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$9221 \$153 \$8115 \$8335 \$8408 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$9224 \$16 \$8436 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9225 \$16 \$8335 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9226 \$16 \$8387 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9227 \$16 \$6989 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9228 \$153 \$8409 \$8230 \$6907 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9229 \$153 \$8409 \$6913 \$8208 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9230 \$16 \$6860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9231 \$16 \$6907 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9232 \$16 \$7466 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9233 \$153 \$8437 \$6719 \$8208 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9234 \$16 \$6979 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9236 \$16 \$8361 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9238 \$16 \$7335 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9240 \$153 \$8362 \$8272 \$6981 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9241 \$153 \$8485 \$6732 \$8363 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9242 \$153 \$8606 \$6913 \$8363 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9244 \$16 \$7992 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9245 \$16 \$7992 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9246 \$16 \$6784 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9247 \$153 \$8439 \$6794 \$8363 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9248 \$16 \$7992 \$16 \$153 \$8363 VNB sky130_fd_sc_hd__inv_1
X$9249 \$16 \$7041 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9252 \$153 \$8458 \$8274 \$7041 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9253 \$16 \$6792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9254 \$153 \$8459 \$8274 \$6860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9255 \$16 \$8364 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9256 \$16 \$7945 \$7887 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$9257 \$153 \$8440 \$6794 \$8196 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9258 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9259 \$16 \$8121 \$7212 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$9260 \$16 \$8121 \$7165 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$9262 \$16 \$8121 \$7156 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$9263 \$16 \$8121 \$8365 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$9264 \$16 \$8422 \$8297 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$9265 \$16 \$8422 \$7655 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$9266 \$16 \$8422 \$8193 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$9267 \$16 \$8340 \$16 \$153 \$8275 VNB sky130_fd_sc_hd__clkbuf_2
X$9268 \$16 \$8275 \$16 \$153 \$8422 VNB sky130_fd_sc_hd__clkbuf_2
X$9269 \$16 \$8275 \$16 \$153 \$8410 VNB sky130_fd_sc_hd__clkbuf_2
X$9270 \$16 \$8422 \$7884 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$9271 \$16 \$8422 \$8335 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$9272 \$16 \$8422 \$8438 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$9273 \$16 \$8212 \$16 \$153 \$8423 VNB sky130_fd_sc_hd__clkbuf_2
X$9274 \$153 \$8411 \$8340 \$6930 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9276 \$153 \$8356 \$8193 \$8386 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$9277 \$16 \$8410 \$6813 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$9279 \$153 \$8460 \$8356 \$6754 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9280 \$16 \$6754 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9281 \$16 \$6930 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9282 \$16 \$6995 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9283 \$153 \$8461 \$8356 \$7044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9285 \$153 \$8442 \$6867 \$8214 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9286 \$16 \$8139 \$7968 \$8462 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$9287 \$153 \$8368 \$8147 \$6916 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9288 \$16 \$8139 \$16 \$153 \$8107 VNB sky130_fd_sc_hd__inv_1
X$9289 \$16 \$6916 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9290 \$153 \$8370 \$8147 \$6771 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9291 \$16 \$8271 \$7968 \$8443 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$9293 \$153 \$7947 \$8335 \$8443 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$9294 \$16 \$8423 \$7968 \$8463 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$9295 \$153 \$8412 \$7947 \$7060 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9296 \$153 \$8388 \$6867 \$8040 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9297 \$153 \$8412 \$6324 \$8040 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9298 \$16 \$8423 \$16 \$153 \$8217 VNB sky130_fd_sc_hd__inv_1
X$9300 \$16 \$8423 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9301 \$16 \$7335 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9302 \$153 \$8464 \$7335 \$8307 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$9303 \$153 \$8279 \$8117 \$8008 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$9304 \$153 \$8444 \$7006 \$8217 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9305 \$153 \$8465 \$8818 \$8424 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9306 \$16 \$7044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9307 \$16 \$7000 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9308 \$16 \$7973 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9310 \$153 \$8413 \$8279 \$6754 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9311 \$153 \$8413 \$6756 \$8218 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9312 \$153 \$8445 \$6324 \$8218 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9313 \$153 \$8466 \$8309 \$6771 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9314 \$16 \$6910 \$8357 \$8414 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$9317 \$16 \$6771 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9318 \$16 \$6910 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9320 \$153 \$8415 \$8309 \$6916 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9321 \$153 \$8390 \$6992 \$8260 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9322 \$153 \$8416 \$6916 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$9323 \$16 \$8416 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9324 \$16 \$6324 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9325 \$16 \$6756 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9327 \$153 \$8415 \$6867 \$8260 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9328 \$153 \$8347 \$6797 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$9329 \$153 \$8467 \$8340 \$6756 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9330 \$16 \$7934 \$7829 \$7949 \$153 \$8078 \$16 VNB sky130_fd_sc_hd__and3b_4
X$9333 \$16 \$7949 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9334 \$153 \$8446 \$8425 \$7067 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9335 \$16 \$7445 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9336 \$16 \$7067 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9338 \$16 \$7328 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9339 \$153 \$8468 \$8425 \$7328 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9340 \$153 \$8446 \$6582 \$8538 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9341 \$16 \$8187 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9342 \$16 \$8673 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9343 \$16 \$7445 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9345 \$153 \$8372 \$8426 \$7445 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9346 \$153 \$8374 \$8426 \$7029 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9347 \$153 \$8375 \$8183 \$7445 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9348 \$16 \$7445 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9349 \$16 \$7029 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9350 \$16 \$8469 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9351 \$16 \$8592 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9353 \$16 \$7239 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9354 \$153 \$8470 \$8183 \$7239 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9356 \$153 \$8183 \$8627 \$8395 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$9358 \$16 \$7029 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9359 \$153 \$8282 \$8281 \$7029 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9360 \$16 \$8731 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9361 \$16 \$7904 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9363 \$153 \$8427 \$7327 \$8263 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9364 \$16 \$8627 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9365 \$16 \$7996 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9366 \$16 \$8819 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9367 \$16 \$7328 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9368 \$153 \$8284 \$8029 \$7328 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9369 \$16 \$7067 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9370 \$16 \$8657 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9372 \$16 \$7029 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9373 \$153 \$8471 \$8184 \$7029 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9375 \$16 \$8624 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9376 \$16 \$7387 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9377 \$153 \$8507 \$8184 \$7387 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9378 \$16 \$8428 \$16 \$153 \$8047 VNB sky130_fd_sc_hd__inv_1
X$9380 \$16 \$7129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9381 \$153 \$8286 \$8030 \$7129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9382 \$16 \$8666 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9383 \$153 \$8076 \$7065 \$8264 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9385 \$16 \$7067 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9387 \$153 \$8472 \$8358 \$7067 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9389 \$16 \$7387 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9390 \$153 \$8474 \$8358 \$7387 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9391 \$16 \$8165 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9392 \$16 \$8165 \$16 \$153 \$8527 VNB sky130_fd_sc_hd__inv_1
X$9393 \$153 \$8030 \$8473 \$8398 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$9394 \$16 \$8165 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9397 \$16 \$8347 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9398 \$16 \$8399 \$16 \$153 \$8165 VNB sky130_fd_sc_hd__clkbuf_2
X$9399 \$153 \$8447 \$8288 \$8245 \$8319 \$8318 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$9400 \$16 \$8049 \$16 \$153 \$8319 VNB sky130_fd_sc_hd__clkbuf_2
X$9401 \$16 \$8050 \$16 \$153 \$8288 VNB sky130_fd_sc_hd__clkbuf_2
X$9402 \$153 \$8347 \$7133 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$9403 \$16 \$8289 \$16 \$153 \$8246 VNB sky130_fd_sc_hd__clkbuf_2
X$9404 \$16 \$8401 \$16 \$153 \$8187 VNB sky130_fd_sc_hd__clkbuf_2
X$9405 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9408 \$153 \$8448 \$8321 \$8225 \$8354 \$8246 \$16 \$16 VNB
+ sky130_fd_sc_hd__nor4b_2
X$9409 \$16 \$8323 \$16 \$153 \$7904 VNB sky130_fd_sc_hd__clkbuf_2
X$9410 \$153 \$8344 \$7208 \$8429 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9411 \$153 \$10311 \$7174 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$9412 \$16 \$7131 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9413 \$153 \$8449 \$7376 \$8378 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9415 \$16 \$7147 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9416 \$153 \$8417 \$8355 \$7147 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9417 \$153 \$8417 \$7463 \$8378 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9419 \$153 \$8418 \$8450 \$7147 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9420 \$153 \$8418 \$7463 \$8380 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9422 \$16 \$7174 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9424 \$153 \$8475 \$8450 \$7174 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9426 \$153 \$8267 \$8290 \$7353 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9427 \$16 \$8044 \$8199 \$8251 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$9429 \$153 \$8476 \$8290 \$7174 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9432 \$16 \$7147 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9433 \$153 \$8477 \$8451 \$7147 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9435 \$16 \$7133 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9436 \$16 \$8165 \$8032 \$8452 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$9437 \$153 \$8031 \$8705 \$8452 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$9438 \$153 \$8478 \$8031 \$7307 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9440 \$16 \$8165 \$16 \$153 \$8291 VNB sky130_fd_sc_hd__inv_1
X$9441 \$153 \$7425 \$7375 \$6985 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9442 \$153 \$7512 \$7462 \$6985 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9443 \$16 \$6985 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9444 \$153 \$8200 \$8732 \$8454 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$9445 \$16 \$8032 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9446 \$16 \$8732 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9448 \$16 \$8453 \$16 \$153 \$8576 VNB sky130_fd_sc_hd__inv_1
X$9449 \$153 \$8430 \$7462 \$8419 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9450 \$16 \$7464 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9452 \$153 \$8420 \$8200 \$7464 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9453 \$153 \$8404 \$7639 \$8291 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9455 \$16 \$7353 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9456 \$16 \$7174 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9457 \$153 \$8479 \$8531 \$7174 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9458 \$153 \$8166 \$7463 \$8576 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9462 \$153 \$8480 \$8330 \$7133 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9463 \$16 \$8704 \$16 \$153 \$8266 VNB sky130_fd_sc_hd__inv_1
X$9464 \$153 \$7517 \$7463 \$7763 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9466 \$16 \$7464 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9467 \$153 \$8455 \$8330 \$7464 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9468 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$9470 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$9471 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$9472 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$9473 \$153 \$8431 \$8331 \$6783 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9474 \$153 \$8510 \$6996 \$8384 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9477 \$16 \$6783 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9479 \$153 \$8532 \$8331 \$6860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9480 \$16 \$6860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9481 \$153 \$8432 \$8331 \$6792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9482 \$16 \$8139 \$16 \$153 \$8384 VNB sky130_fd_sc_hd__inv_1
X$9483 \$153 \$8481 \$8333 \$6907 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9485 \$16 \$6907 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9487 \$153 \$8511 \$6996 \$8206 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9488 \$153 \$8482 \$8333 \$6784 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9489 \$153 \$8333 \$8503 \$8421 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$9490 \$153 \$8533 \$7659 \$8633 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$9492 \$16 \$7521 \$16 \$153 \$8723 VNB sky130_fd_sc_hd__inv_1
X$9493 \$16 \$6784 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9495 \$153 \$8535 \$8387 \$8534 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$9496 \$153 \$8483 \$8457 \$8723 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9497 \$16 \$8580 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9498 \$153 \$8484 \$8230 \$7041 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9499 \$153 \$8484 \$6996 \$8208 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9501 \$153 \$8437 \$8230 \$6792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9502 \$16 \$7466 \$8504 \$8536 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$9503 \$16 \$6792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9504 \$153 \$8485 \$8272 \$6860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9505 \$16 \$6783 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9506 \$16 \$6860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9508 \$16 \$6981 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9509 \$153 \$8512 \$8457 \$8513 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9512 \$153 \$8486 \$8272 \$7041 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9513 \$153 \$8486 \$6996 \$8363 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9514 \$153 \$8211 \$8274 \$6907 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9515 \$16 \$6907 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9517 \$153 \$8514 \$8737 \$8515 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9518 \$16 \$8177 \$16 \$153 \$8196 VNB sky130_fd_sc_hd__inv_1
X$9520 \$153 \$8458 \$6996 \$8196 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9521 \$16 \$8410 \$7333 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$9522 \$153 \$8301 \$6783 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$9523 \$153 \$8516 \$6981 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$9524 \$16 \$8422 \$8167 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$9527 \$16 \$8410 \$7237 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$9528 \$16 \$8410 \$6888 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$9529 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9530 \$153 \$8441 \$8340 \$6719 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9531 \$153 \$8487 \$8340 \$6995 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9532 \$153 \$8367 \$8356 \$6797 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9534 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9535 \$16 \$6797 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9536 \$153 \$8460 \$6756 \$8214 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9538 \$153 \$8442 \$8356 \$6916 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9539 \$153 \$8461 \$7006 \$8214 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9540 \$16 \$6916 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9542 \$153 \$8147 \$8167 \$8462 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$9544 \$16 \$8139 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9546 \$16 \$8387 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9547 \$16 \$8635 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9548 \$153 \$8369 \$8147 \$7044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9549 \$153 \$8587 \$8387 \$8517 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$9550 \$16 \$7521 \$8635 \$8518 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$9551 \$153 \$8278 \$8503 \$8463 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$9553 \$16 \$8503 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9555 \$153 \$8488 \$8278 \$6771 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9556 \$153 \$8488 \$6865 \$8217 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9557 \$16 \$6771 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9558 \$153 \$8505 \$6756 \$8217 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9559 \$153 \$8537 \$8278 \$7060 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9562 \$16 \$7060 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9564 \$153 \$8371 \$8279 \$6771 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9565 \$16 \$7000 \$8357 \$8519 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$9566 \$16 \$6771 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9568 \$153 \$8489 \$8279 \$6797 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9569 \$153 \$8489 \$6906 \$8218 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9570 \$16 \$6754 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9571 \$16 \$6797 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9573 \$16 \$7000 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9574 \$16 \$7226 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9575 \$153 \$7898 \$8309 \$7044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9576 \$153 \$8466 \$6865 \$8260 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9577 \$16 \$7044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9578 \$16 \$6935 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9579 \$153 \$8490 \$8309 \$7060 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9580 \$16 \$6916 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9581 \$16 \$7060 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9582 \$16 \$8686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9585 \$153 \$8520 \$8610 \$8613 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9586 \$16 \$8556 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9587 \$153 \$8734 \$7060 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$9588 \$153 \$10383 \$7044 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$9589 \$16 \$10383 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9591 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9593 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9594 \$153 \$8521 \$9278 \$7994 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9595 \$153 \$8491 \$8340 \$6992 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9596 \$16 \$6906 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9597 \$153 \$8492 \$8425 \$7445 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9598 \$153 \$8392 \$6582 \$7860 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9599 \$16 \$7029 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9601 \$153 \$8493 \$8425 \$7029 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9602 \$16 \$7129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9603 \$16 \$7239 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9604 \$153 \$8494 \$8426 \$7129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9605 \$153 \$8493 \$7066 \$8538 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9606 \$153 \$8522 \$7482 \$8373 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9607 \$16 \$8539 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9610 \$153 \$8495 \$8183 \$7029 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9612 \$16 \$8523 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9613 \$16 \$8540 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9614 \$16 \$8524 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9615 \$153 \$8620 \$4675 \$8341 \$8523 \$7834 \$8506 \$8593 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$9616 \$16 \$8541 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9617 \$153 \$8394 \$7490 \$8043 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9619 \$16 \$7996 \$16 \$153 \$8043 VNB sky130_fd_sc_hd__inv_1
X$9620 \$153 \$7997 \$7215 \$8222 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9621 \$153 \$8542 \$8281 \$7328 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9622 \$16 \$7328 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9623 \$16 \$7239 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9624 \$153 \$8376 \$8029 \$7239 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9625 \$16 \$7130 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9626 \$16 \$7130 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9627 \$16 \$7994 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9628 \$16 \$7994 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9630 \$153 \$8752 \$7215 \$8525 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9631 \$16 \$8316 \$16 \$153 \$8222 VNB sky130_fd_sc_hd__inv_1
X$9632 \$153 \$8029 \$8285 \$8526 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$9633 \$153 \$8349 \$8184 \$7067 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9634 \$16 \$8624 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9636 \$153 \$8507 \$7490 \$8047 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9637 \$16 \$8428 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9639 \$153 \$8184 \$8666 \$8543 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$9640 \$16 \$7328 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9641 \$153 \$8496 \$8358 \$7328 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9643 \$153 \$8496 \$7366 \$8527 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9644 \$153 \$8472 \$6582 \$8527 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9646 \$16 \$8473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9647 \$16 \$8198 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9650 \$16 \$8359 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9651 \$16 \$7239 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9652 \$153 \$8474 \$7490 \$8527 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9653 \$153 \$8497 \$7482 \$8527 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9655 \$16 \$8287 \$16 \$153 \$8265 VNB sky130_fd_sc_hd__clkbuf_2
X$9656 \$16 \$8447 \$16 \$153 \$8704 VNB sky130_fd_sc_hd__clkbuf_2
X$9657 \$16 \$8528 \$16 \$153 \$8453 VNB sky130_fd_sc_hd__clkbuf_2
X$9658 \$153 \$8544 \$8318 \$8319 \$8288 \$8245 \$16 \$16 VNB
+ sky130_fd_sc_hd__nor4b_2
X$9659 \$16 \$8245 \$8288 \$8319 \$8318 \$16 \$153 \$8545 VNB
+ sky130_fd_sc_hd__and4_2
X$9661 \$153 \$8320 \$7147 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$9662 \$153 \$8546 \$8225 \$8246 \$8321 \$8354 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$9663 \$153 \$8547 \$8354 \$8246 \$8225 \$8321 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$9664 \$153 \$8506 \$8340 \$7208 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9666 \$16 \$10311 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9667 \$16 \$7463 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9669 \$16 \$7377 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9670 \$153 \$8449 \$8355 \$7174 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9671 \$16 \$7174 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9672 \$16 \$7376 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9674 \$16 \$7133 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9675 \$153 \$8499 \$8355 \$7133 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9676 \$153 \$8499 \$7180 \$8378 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9679 \$153 \$8379 \$8450 \$7133 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9680 \$16 \$7133 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9681 \$16 \$7307 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9682 \$153 \$8381 \$8450 \$7131 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9683 \$153 \$8475 \$7376 \$8380 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9684 \$16 \$7147 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9685 \$153 \$8383 \$7375 \$8266 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9687 \$153 \$8500 \$8290 \$7147 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9688 \$153 \$8500 \$7463 \$8268 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9689 \$16 \$7174 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9691 \$16 \$7174 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9692 \$153 \$8549 \$8451 \$7174 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9693 \$153 \$8477 \$7463 \$8529 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9696 \$153 \$8501 \$8451 \$7133 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9697 \$153 \$8501 \$7180 \$8529 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9699 \$16 \$7147 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9700 \$153 \$8502 \$8508 \$7131 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9701 \$153 \$8502 \$7208 \$8419 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9703 \$16 \$7133 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9705 \$16 \$8453 \$8032 \$8454 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$9707 \$153 \$8550 \$8508 \$7133 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9708 \$153 \$8530 \$7376 \$8419 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9709 \$16 \$8351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9710 \$16 \$8353 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9711 \$16 \$7147 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9712 \$153 \$8498 \$8531 \$7147 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9714 \$16 \$7131 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9717 \$153 \$8344 \$8531 \$7131 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9718 \$153 \$8330 \$8353 \$8509 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$9719 \$16 \$8704 \$8032 \$8509 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$9720 \$153 \$7843 \$7208 \$7763 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9721 \$153 \$7682 \$7375 \$7763 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9722 \$16 \$7131 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9724 \$16 \$8704 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9726 \$16 \$7377 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9727 \$153 \$8551 \$8330 \$7377 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9728 \$153 \$7764 \$7639 \$7763 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9729 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$9730 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$9732 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$9733 \$153 \$11048 \$10962 \$10295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9734 \$153 \$10997 \$10327 \$11055 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9735 \$16 \$10295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9736 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$9737 \$153 \$11071 \$10962 \$10367 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9738 \$16 \$10367 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9739 \$16 \$10646 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9740 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$9742 \$153 \$11071 \$10330 \$11055 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9743 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$9744 \$16 \$10476 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9745 \$153 \$10962 \$11004 \$11072 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$9746 \$16 \$11004 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9747 \$16 \$11078 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9749 \$153 \$10964 \$10963 \$10226 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9750 \$16 \$10226 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9751 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$9753 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$9754 \$153 \$10965 \$10963 \$10367 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9756 \$153 \$11073 \$10303 \$10884 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9758 \$153 \$10532 \$11114 \$10998 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$9760 \$153 \$11074 \$10088 \$10745 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9764 \$153 \$10967 \$10966 \$10226 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9765 \$16 \$10646 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9767 \$153 \$11075 \$10966 \$10368 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9768 \$153 \$11075 \$10303 \$11056 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9769 \$16 \$10368 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9770 \$153 \$11076 \$10705 \$11056 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9772 \$16 \$11077 \$10635 \$11115 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$9773 \$16 \$11077 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9775 \$153 \$11116 \$11000 \$10368 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9776 \$16 \$10368 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9777 \$153 \$10969 \$11000 \$10295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9778 \$153 \$11116 \$10303 \$10954 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9779 \$16 \$10295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9780 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$9782 \$153 \$11179 \$10971 \$10646 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9783 \$153 \$11117 \$10971 \$10295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9784 \$153 \$11117 \$10276 \$11057 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9785 \$16 \$10295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9786 \$16 \$11267 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9787 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$9789 \$16 \$10974 \$16 \$153 \$10805 VNB sky130_fd_sc_hd__inv_1
X$9793 \$16 \$11118 \$16 \$153 \$11077 VNB sky130_fd_sc_hd__clkbuf_2
X$9794 \$16 \$10974 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9795 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$9797 \$153 \$11003 \$10088 \$10805 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9798 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$9799 \$16 \$11111 \$16 \$153 \$10907 VNB sky130_fd_sc_hd__clkbuf_2
X$9800 \$153 \$11058 \$10907 \$10878 \$10877 \$10885 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$9801 \$16 \$10878 \$10907 \$10877 \$10885 \$16 \$153 \$11136 VNB
+ sky130_fd_sc_hd__and4_2
X$9802 \$16 \$6667 \$16 \$153 \$11119 VNB sky130_fd_sc_hd__clkbuf_2
X$9803 \$16 \$11079 \$16 \$153 \$10939 VNB sky130_fd_sc_hd__clkbuf_2
X$9806 \$16 \$11078 \$10525 \$11080 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$9807 \$16 \$11078 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9808 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$9810 \$153 \$11137 \$11120 \$10606 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9811 \$16 \$10606 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9812 \$153 \$11081 \$10686 \$10941 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9813 \$16 \$10605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9815 \$16 \$10764 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9816 \$153 \$11082 \$10309 \$10941 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9817 \$16 \$10338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9820 \$153 \$11059 \$10821 \$10470 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9821 \$16 \$10298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9822 \$16 \$10382 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9824 \$153 \$11138 \$11121 \$10382 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9826 \$153 \$11122 \$10401 \$11112 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9827 \$153 \$11005 \$10538 \$10750 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9829 \$16 \$10939 \$10525 \$11083 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$9830 \$16 \$11123 \$16 \$153 \$10525 VNB sky130_fd_sc_hd__clkbuf_2
X$9831 \$16 \$10514 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9832 \$153 \$10972 \$11060 \$10470 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9833 \$16 \$10939 \$16 \$153 \$10956 VNB sky130_fd_sc_hd__inv_1
X$9834 \$16 \$10470 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9835 \$16 \$10939 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9837 \$153 \$10973 \$11060 \$10382 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9839 \$16 \$10514 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9840 \$16 \$10382 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9843 \$16 \$11123 \$16 \$153 \$10655 VNB sky130_fd_sc_hd__clkbuf_2
X$9844 \$153 \$11139 \$11124 \$10470 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9845 \$153 \$11036 \$10344 \$10958 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9846 \$16 \$10470 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9847 \$153 \$10957 \$11124 \$10298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9848 \$16 \$10338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9849 \$16 \$10298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9850 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$9852 \$153 \$11140 \$11049 \$10526 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9853 \$16 \$10526 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9854 \$16 \$11488 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9856 \$153 \$11084 \$11049 \$10605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9857 \$153 \$11125 \$10401 \$11061 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9858 \$153 \$11084 \$10686 \$11061 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9861 \$153 \$11141 \$10893 \$10514 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9862 \$153 \$11086 \$10893 \$10606 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9863 \$153 \$11086 \$10344 \$10892 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9864 \$153 \$11085 \$10686 \$10892 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9865 \$16 \$10606 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9867 \$16 \$10974 \$16 \$153 \$10894 VNB sky130_fd_sc_hd__inv_1
X$9869 \$153 \$11087 \$10401 \$10894 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9870 \$153 \$11126 \$10344 \$10894 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9872 \$153 \$11063 \$10975 \$10526 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9873 \$153 \$11142 \$10975 \$10605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9874 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$9875 \$16 \$10473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9877 \$153 \$11064 \$11050 \$10473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9879 \$16 \$10611 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9880 \$16 \$10386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9881 \$16 \$10809 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9882 \$153 \$11143 \$11050 \$10386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9883 \$153 \$11144 \$10734 \$10809 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9885 \$153 \$11128 \$10370 \$11207 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9886 \$16 \$10551 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9887 \$153 \$10977 \$10734 \$10551 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9888 \$16 \$10978 \$11127 \$11145 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$9889 \$153 \$11146 \$10979 \$10809 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9890 \$16 \$10978 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9891 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$9894 \$16 \$10300 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9895 \$153 \$11092 \$10979 \$10300 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9896 \$153 \$11092 \$10417 \$10810 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9897 \$16 \$9200 \$16 \$153 \$11212 VNB sky130_fd_sc_hd__clkbuf_2
X$9899 \$153 \$11093 \$10881 \$10578 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9900 \$16 \$10578 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9901 \$16 \$10809 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9902 \$16 \$11214 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9904 \$153 \$11093 \$10370 \$10946 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9905 \$16 \$10611 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9906 \$16 \$10551 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9907 \$153 \$11094 \$10882 \$10551 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9908 \$153 \$11129 \$10882 \$10809 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9909 \$153 \$11129 \$10714 \$10811 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9910 \$16 \$10300 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9913 \$153 \$10922 \$10501 \$10811 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9915 \$16 \$10809 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9916 \$153 \$11095 \$10834 \$10809 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9918 \$153 \$11095 \$10714 \$10923 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9919 \$153 \$11130 \$10501 \$10948 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9920 \$16 \$10551 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9921 \$16 \$12050 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9922 \$16 \$10649 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9923 \$16 \$10735 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9925 \$153 \$10984 \$10834 \$10735 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9926 \$16 \$10386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9927 \$153 \$11131 \$10833 \$11099 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9928 \$153 \$11132 \$11066 \$10386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9929 \$153 \$10692 \$10833 \$10926 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9931 \$16 \$11172 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9934 \$16 \$10300 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9935 \$16 \$11172 \$16 \$153 \$11099 VNB sky130_fd_sc_hd__inv_1
X$9936 \$153 \$11097 \$11066 \$10300 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9938 \$153 \$11098 \$10714 \$11099 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9939 \$153 \$11097 \$10417 \$11099 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9940 \$16 \$6667 \$16 \$153 \$11147 VNB sky130_fd_sc_hd__clkbuf_2
X$9941 \$16 \$11133 \$16 \$153 \$11113 VNB sky130_fd_sc_hd__clkbuf_2
X$9942 \$16 \$11188 \$16 \$153 \$10978 VNB sky130_fd_sc_hd__clkbuf_2
X$9943 \$16 \$6667 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9947 \$16 \$11113 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9948 \$153 \$11012 \$10987 \$10929 \$10950 \$10988 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$9949 \$16 \$10988 \$10987 \$11012 \$10950 \$16 \$153 \$11069 VNB
+ sky130_fd_sc_hd__and4_2
X$9950 \$16 \$11148 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9951 \$153 \$11102 \$10466 \$11016 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9952 \$153 \$11014 \$10815 \$10812 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9953 \$153 \$11149 \$11052 \$10392 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9955 \$16 \$10978 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9956 \$16 \$11016 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9958 \$153 \$11134 \$10642 \$10961 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9960 \$153 \$11101 \$11052 \$10467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9961 \$16 \$10467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9962 \$16 \$11102 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9964 \$16 \$12347 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9965 \$153 \$11103 \$11052 \$10393 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9966 \$16 \$10393 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9968 \$153 \$11103 \$10694 \$10961 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9969 \$16 \$11013 \$16 \$153 \$10814 VNB sky130_fd_sc_hd__inv_1
X$9970 \$153 \$10991 \$10740 \$10617 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9971 \$16 \$10617 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9973 \$153 \$10993 \$10740 \$10467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9974 \$153 \$11104 \$10642 \$10814 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9976 \$153 \$11150 \$10901 \$10446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9977 \$16 \$10446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9978 \$16 \$10467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9979 \$153 \$11151 \$10901 \$10467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9981 \$153 \$10995 \$10615 \$11018 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$9982 \$16 \$10615 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9984 \$16 \$10649 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9986 \$16 \$10552 \$16 \$153 \$11516 VNB sky130_fd_sc_hd__inv_1
X$9987 \$153 \$10934 \$10587 \$10858 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9988 \$153 \$10420 \$10285 \$10858 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9989 \$153 \$10628 \$10642 \$10858 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$9991 \$16 \$10392 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9992 \$153 \$11152 \$10995 \$10392 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$9993 \$16 \$10853 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9995 \$16 \$10960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9996 \$16 \$10392 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$9998 \$153 \$10448 \$10376 \$10650 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10000 \$16 \$10393 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10002 \$16 \$10446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10003 \$153 \$11153 \$11053 \$10446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10004 \$16 \$10222 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10006 \$16 \$10326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10007 \$16 \$10346 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10009 \$153 \$11135 \$11053 \$10326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10012 \$153 \$10800 \$10694 \$10741 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10013 \$153 \$10799 \$10285 \$10741 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10015 \$16 \$10392 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10016 \$153 \$10633 \$10376 \$10741 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10017 \$153 \$11154 \$10796 \$10392 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10019 \$153 \$9992 \$9103 \$10510 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10021 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$10022 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$10023 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$10025 \$153 \$11231 \$11288 \$10295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10026 \$16 \$10295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10027 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$10029 \$153 \$11155 \$10962 \$10646 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10030 \$153 \$11155 \$10318 \$11055 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10031 \$153 \$11189 \$10330 \$11232 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10032 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$10033 \$153 \$11176 \$10161 \$11232 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10036 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$10038 \$153 \$11234 \$10963 \$10476 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10039 \$16 \$10368 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10040 \$16 \$10476 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10042 \$16 \$10427 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10043 \$153 \$11156 \$10963 \$10427 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10044 \$16 \$10367 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10046 \$16 \$11274 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10047 \$16 \$10200 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10049 \$153 \$11156 \$10327 \$10884 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10050 \$16 \$11274 \$11347 \$11236 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$10052 \$16 \$11190 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10053 \$16 \$11274 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10054 \$16 \$11114 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10056 \$153 \$11192 \$10276 \$11191 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10057 \$153 \$11193 \$10303 \$11191 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10058 \$153 \$11157 \$10966 \$10200 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10061 \$153 \$11157 \$10088 \$11056 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10062 \$153 \$11177 \$10276 \$11393 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10063 \$16 \$11077 \$16 \$153 \$11056 VNB sky130_fd_sc_hd__inv_1
X$10064 \$153 \$10966 \$11194 \$11115 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$10065 \$16 \$10953 \$16 \$153 \$10635 VNB sky130_fd_sc_hd__clkbuf_2
X$10066 \$16 \$10953 \$16 \$153 \$11238 VNB sky130_fd_sc_hd__clkbuf_2
X$10067 \$16 \$11194 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10068 \$16 \$11077 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10069 \$16 \$9200 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10070 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$10072 \$153 \$11239 \$10327 \$10954 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10073 \$16 \$11240 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10075 \$153 \$11178 \$10088 \$10954 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10076 \$153 \$11158 \$10971 \$10226 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10078 \$153 \$11179 \$10318 \$11057 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10079 \$16 \$10646 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10080 \$16 \$10226 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10081 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$10083 \$153 \$11195 \$10327 \$11057 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10084 \$16 \$11267 \$16 \$153 \$11057 VNB sky130_fd_sc_hd__inv_1
X$10085 \$16 \$10200 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10086 \$153 \$10817 \$10959 \$11242 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$10087 \$16 \$10959 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10088 \$153 \$11196 \$11243 \$11159 \$11197 \$11180 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$10089 \$153 \$11181 \$10276 \$10805 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10090 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$10092 \$16 \$6540 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10095 \$16 \$11119 \$16 \$153 \$10885 VNB sky130_fd_sc_hd__clkbuf_2
X$10097 \$16 \$6540 \$16 \$153 \$11111 VNB sky130_fd_sc_hd__clkbuf_2
X$10098 \$16 \$7559 \$16 \$153 \$11244 VNB sky130_fd_sc_hd__clkbuf_2
X$10099 \$16 \$11244 \$16 \$153 \$10877 VNB sky130_fd_sc_hd__clkbuf_2
X$10101 \$16 \$11198 \$16 \$153 \$10878 VNB sky130_fd_sc_hd__clkbuf_2
X$10102 \$16 \$11136 \$16 \$153 \$10730 VNB sky130_fd_sc_hd__clkbuf_2
X$10103 \$16 \$11199 \$16 \$153 \$11159 VNB sky130_fd_sc_hd__clkbuf_2
X$10104 \$16 \$7559 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10105 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$10106 \$16 \$7656 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10108 \$153 \$11160 \$11120 \$10526 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10112 \$153 \$11160 \$10516 \$11200 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10113 \$153 \$11298 \$10538 \$11200 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10114 \$153 \$11161 \$11120 \$10298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10115 \$153 \$11161 \$10401 \$11200 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10116 \$153 \$11182 \$10098 \$11200 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10117 \$16 \$10298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10120 \$153 \$11245 \$11121 \$10338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10121 \$16 \$10338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10123 \$16 \$10744 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10124 \$153 \$11162 \$11121 \$10514 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10125 \$153 \$11162 \$10538 \$11112 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10127 \$153 \$11201 \$10344 \$10956 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10129 \$16 \$10526 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10131 \$16 \$10338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10133 \$153 \$11163 \$11060 \$10514 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10134 \$153 \$11163 \$10538 \$10956 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10135 \$153 \$11183 \$10686 \$10956 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10136 \$16 \$11123 \$16 \$153 \$11164 VNB sky130_fd_sc_hd__clkbuf_2
X$10138 \$153 \$11202 \$10538 \$10958 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10140 \$153 \$11184 \$10516 \$10958 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10141 \$153 \$11139 \$10247 \$10958 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10142 \$153 \$11203 \$10686 \$10958 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10143 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$10144 \$153 \$11204 \$10247 \$11488 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10145 \$153 \$11140 \$10516 \$11061 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10146 \$16 \$10338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10147 \$16 \$11077 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10148 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$10150 \$153 \$11125 \$11049 \$10298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10151 \$16 \$10298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10152 \$153 \$11062 \$10893 \$10338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10154 \$153 \$11141 \$10538 \$10892 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10155 \$153 \$11247 \$10247 \$11205 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10156 \$16 \$10514 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10159 \$153 \$10975 \$10959 \$11206 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$10160 \$153 \$11126 \$10975 \$10606 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10162 \$153 \$11165 \$10501 \$11207 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10163 \$153 \$11248 \$11208 \$10605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10165 \$16 \$11207 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10167 \$153 \$11248 \$10686 \$11268 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10168 \$16 \$10605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10170 \$16 \$10300 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10171 \$153 \$11166 \$11050 \$10300 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10173 \$153 \$11088 \$10714 \$11209 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10174 \$153 \$11166 \$10417 \$11209 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10175 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$10177 \$153 \$11210 \$10370 \$11209 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10178 \$153 \$11143 \$10472 \$11209 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10179 \$16 \$11113 \$11127 \$11250 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$10181 \$153 \$11090 \$11185 \$10386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10183 \$153 \$10734 \$11015 \$11145 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$10186 \$16 \$10611 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10187 \$16 \$10551 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10188 \$153 \$10832 \$10979 \$10611 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10189 \$153 \$11144 \$10714 \$10480 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10190 \$153 \$11211 \$10471 \$10810 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10191 \$153 \$11009 \$10472 \$10810 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10192 \$16 \$11212 \$16 \$153 \$11127 VNB sky130_fd_sc_hd__clkbuf_2
X$10193 \$16 \$10300 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10194 \$16 \$11013 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10196 \$16 \$9200 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10197 \$16 \$10473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10198 \$153 \$11213 \$10472 \$10946 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10199 \$153 \$11186 \$10714 \$10946 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10200 \$153 \$11186 \$10881 \$10809 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10201 \$16 \$11214 \$16 \$153 \$10946 VNB sky130_fd_sc_hd__inv_1
X$10202 \$153 \$11333 \$10833 \$11215 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10203 \$16 \$11216 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10204 \$16 \$11214 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10207 \$16 \$10809 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10208 \$16 \$10578 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10209 \$153 \$11167 \$10882 \$10578 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10210 \$153 \$11167 \$10370 \$10811 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10211 \$153 \$10559 \$10417 \$10757 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10212 \$153 \$10503 \$10501 \$10757 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10213 \$153 \$10690 \$10833 \$10757 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10215 \$153 \$11217 \$10714 \$10948 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10216 \$16 \$10649 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10217 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$10218 \$153 \$11218 \$10471 \$11219 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10219 \$153 \$11187 \$10919 \$11219 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10220 \$153 \$11220 \$10501 \$11219 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10222 \$16 \$10473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10223 \$153 \$11168 \$10501 \$11099 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10225 \$153 \$11168 \$11066 \$10473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10226 \$153 \$11096 \$10370 \$11099 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10227 \$153 \$11132 \$10472 \$11099 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10228 \$16 \$10551 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10229 \$153 \$11169 \$11066 \$10551 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10230 \$16 \$11221 \$16 \$153 \$10988 VNB sky130_fd_sc_hd__clkbuf_2
X$10232 \$153 \$11169 \$10471 \$11099 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10233 \$16 \$7559 \$16 \$153 \$11253 VNB sky130_fd_sc_hd__clkbuf_2
X$10234 \$16 \$11147 \$16 \$153 \$11222 VNB sky130_fd_sc_hd__clkbuf_2
X$10235 \$153 \$11188 \$11254 \$11223 \$11255 \$11222 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$10236 \$16 \$11253 \$16 \$153 \$11255 VNB sky130_fd_sc_hd__clkbuf_2
X$10238 \$153 \$11255 \$11254 \$11224 \$11222 \$11223 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$10240 \$16 \$11113 \$10838 \$11170 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$10241 \$153 \$11318 \$10694 \$11016 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10243 \$153 \$11052 \$11148 \$11170 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$10244 \$16 \$10978 \$16 \$153 \$10812 VNB sky130_fd_sc_hd__inv_1
X$10245 \$153 \$11134 \$11052 \$10564 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10246 \$153 \$11225 \$10466 \$11226 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10247 \$153 \$11149 \$10815 \$10961 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10248 \$16 \$11113 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10250 \$16 \$11013 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10252 \$16 \$10446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10253 \$16 \$10393 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10254 \$153 \$11257 \$11052 \$10446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10256 \$153 \$10740 \$12347 \$11258 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$10257 \$153 \$11227 \$10376 \$11384 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10258 \$153 \$10933 \$10815 \$10814 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10260 \$16 \$11216 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10262 \$16 \$10467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10264 \$16 \$10990 \$16 \$153 \$11504 VNB sky130_fd_sc_hd__clkbuf_2
X$10265 \$153 \$10901 \$11216 \$11259 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$10266 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$10267 \$16 \$11214 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10268 \$153 \$11228 \$10466 \$11495 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10269 \$16 \$11214 \$16 \$153 \$10902 VNB sky130_fd_sc_hd__inv_1
X$10270 \$153 \$11150 \$10376 \$10902 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10271 \$153 \$11105 \$10642 \$11516 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10273 \$153 \$11171 \$10901 \$10326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10274 \$153 \$11151 \$10587 \$10902 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10275 \$153 \$11171 \$10466 \$10902 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10276 \$16 \$10552 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10278 \$153 \$10447 \$10376 \$10858 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10279 \$153 \$10697 \$10694 \$10858 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10281 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$10282 \$16 \$11172 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10283 \$16 \$10446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10284 \$153 \$10794 \$10815 \$10650 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10285 \$153 \$11261 \$11285 \$10446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10287 \$16 \$10467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10288 \$16 \$11172 \$11229 \$11262 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$10289 \$153 \$11173 \$11053 \$10467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10291 \$16 \$10529 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10293 \$16 \$10392 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10294 \$16 \$10617 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10296 \$153 \$11174 \$11053 \$10392 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10297 \$153 \$10841 \$10642 \$11022 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10298 \$153 \$11590 \$11230 \$10564 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10299 \$16 \$10564 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10300 \$16 \$11172 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10301 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$10303 \$16 \$10467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10304 \$16 \$10446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10305 \$16 \$10617 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10306 \$153 \$11175 \$11230 \$10617 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10307 \$153 \$10055 \$8965 \$10510 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10308 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$10309 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$10311 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$10312 \$153 \$4967 \$4864 \$3766 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10313 \$153 \$4967 \$3478 \$4859 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10314 \$153 \$5021 \$3394 \$4859 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10315 \$153 \$4469 \$5152 \$5022 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$10316 \$16 \$4742 \$4538 \$5022 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$10318 \$16 \$4538 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10320 \$153 \$5047 \$4788 \$3571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10321 \$153 \$5048 \$4788 \$3385 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10322 \$16 \$4893 \$4538 \$5049 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$10324 \$153 \$4969 \$3478 \$4692 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10325 \$16 \$5080 \$4538 \$5050 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$10328 \$153 \$5048 \$3394 \$4692 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10329 \$153 \$4894 \$3394 \$4707 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10330 \$16 \$5080 \$16 \$153 \$4707 VNB sky130_fd_sc_hd__inv_1
X$10331 \$16 \$4538 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10332 \$16 \$3385 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10333 \$153 \$5052 \$4789 \$3385 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10334 \$153 \$4895 \$3606 \$4693 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10335 \$16 \$3571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10337 \$16 \$4896 \$16 \$153 \$4693 VNB sky130_fd_sc_hd__inv_1
X$10339 \$153 \$4789 \$4939 \$5023 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$10340 \$153 \$4897 \$3540 \$4693 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10342 \$16 \$4947 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10343 \$16 \$3571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10344 \$153 \$4972 \$3606 \$4940 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10345 \$153 \$4813 \$3307 \$4940 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10347 \$153 \$5024 \$3422 \$4359 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10349 \$153 \$4899 \$3540 \$4940 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10350 \$16 \$3616 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10351 \$16 \$4947 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10352 \$16 \$4538 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10353 \$153 \$5053 \$4867 \$3385 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10354 \$16 \$3385 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10356 \$153 \$5054 \$5055 \$5168 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10357 \$153 \$4900 \$3606 \$4359 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10358 \$16 \$5026 \$16 \$153 \$4359 VNB sky130_fd_sc_hd__inv_1
X$10361 \$16 \$5026 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10362 \$16 \$3766 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10363 \$153 \$5056 \$4791 \$3766 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10364 \$153 \$5057 \$4791 \$3385 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10366 \$16 \$4869 \$16 \$153 \$4941 VNB sky130_fd_sc_hd__inv_1
X$10367 \$153 \$4791 \$5228 \$4975 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$10368 \$16 \$3709 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10370 \$16 \$5228 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10371 \$16 \$4869 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10372 \$16 \$3571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10373 \$153 \$5025 \$3422 \$4694 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10374 \$153 \$4944 \$4711 \$3766 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10375 \$16 \$3766 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10377 \$16 \$4976 \$16 \$153 \$5026 VNB sky130_fd_sc_hd__clkbuf_2
X$10378 \$153 \$4659 \$4714 \$5058 \$4715 \$4598 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$10379 \$153 \$4715 \$4714 \$5059 \$4659 \$4598 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$10381 \$16 \$4598 \$4714 \$4659 \$4715 \$16 \$153 \$4946 VNB
+ sky130_fd_sc_hd__and4_2
X$10383 \$16 \$4977 \$16 \$153 \$4947 VNB sky130_fd_sc_hd__clkbuf_2
X$10384 \$153 \$5027 \$4661 \$4662 \$4717 \$4716 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$10385 \$153 \$4599 \$5226 \$5028 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$10386 \$16 \$4742 \$4275 \$5060 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$10387 \$16 \$4275 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10388 \$16 \$4742 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10389 \$16 \$3778 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10391 \$16 \$4742 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10392 \$16 \$4742 \$16 \$153 \$4861 VNB sky130_fd_sc_hd__inv_1
X$10393 \$16 \$4902 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10395 \$16 \$3621 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10396 \$153 \$4979 \$4926 \$3543 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10397 \$153 \$4979 \$3556 \$4861 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10398 \$16 \$3543 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10399 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$10400 \$16 \$5051 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10401 \$153 \$5029 \$3504 \$4861 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10402 \$153 \$5030 \$3354 \$4861 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10404 \$16 \$5080 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10407 \$16 \$5080 \$16 \$153 \$4796 VNB sky130_fd_sc_hd__inv_1
X$10408 \$153 \$5031 \$5209 \$5564 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10409 \$153 \$5032 \$3101 \$4796 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10410 \$153 \$5033 \$5209 \$5013 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10411 \$153 \$5034 \$3504 \$4796 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10412 \$153 \$5061 \$4797 \$3492 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10414 \$16 \$4896 \$16 \$153 \$4818 VNB sky130_fd_sc_hd__inv_1
X$10415 \$153 \$5035 \$3504 \$4818 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10416 \$16 \$3492 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10417 \$16 \$4275 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10418 \$16 \$4893 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10419 \$153 \$5062 \$4797 \$3572 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10420 \$16 \$4893 \$16 \$153 \$4530 VNB sky130_fd_sc_hd__inv_1
X$10421 \$16 \$3621 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10423 \$153 \$5063 \$4622 \$3492 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10425 \$16 \$3492 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10426 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$10427 \$153 \$5036 \$3101 \$4530 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10428 \$153 \$5063 \$3354 \$4530 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10429 \$16 \$3543 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10430 \$153 \$5014 \$3556 \$4798 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10431 \$16 \$4947 \$16 \$153 \$4798 VNB sky130_fd_sc_hd__inv_1
X$10432 \$16 \$4947 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10433 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$10435 \$153 \$4821 \$3354 \$4798 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10436 \$16 \$3572 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10439 \$16 \$5026 \$3957 \$5064 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$10440 \$16 \$5026 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10441 \$16 \$4943 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10442 \$153 \$4981 \$3079 \$4696 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10443 \$153 \$5037 \$3504 \$4696 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10444 \$153 \$4905 \$3354 \$4696 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10445 \$16 \$5026 \$16 \$153 \$4696 VNB sky130_fd_sc_hd__inv_1
X$10447 \$153 \$5038 \$3101 \$4696 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10448 \$16 \$5026 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10449 \$16 \$4712 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10451 \$16 \$5065 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10453 \$16 \$4869 \$3957 \$4824 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$10454 \$16 \$4869 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10455 \$16 \$4822 \$16 \$153 \$5066 VNB sky130_fd_sc_hd__inv_1
X$10456 \$16 \$4822 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10457 \$153 \$4982 \$3608 \$5066 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10458 \$16 \$3572 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10459 \$16 \$3241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10460 \$153 \$5067 \$4948 \$3480 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10462 \$153 \$153 \$5519 \$5155 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10463 \$16 \$4983 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10465 \$16 \$3492 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10467 \$153 \$5068 \$4948 \$3492 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10468 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$10469 \$16 \$5069 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10470 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10471 \$153 \$3674 \$1482 \$5069 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10472 \$153 \$5068 \$3354 \$5066 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10473 \$16 \$4048 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10474 \$16 \$3889 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10476 \$16 \$3731 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10478 \$153 \$4929 \$4799 \$3792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10479 \$153 \$4802 \$4799 \$3814 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10480 \$16 \$4760 \$16 \$153 \$4801 VNB sky130_fd_sc_hd__inv_1
X$10481 \$16 \$5452 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10483 \$153 \$4985 \$3763 \$4801 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10484 \$153 \$4986 \$3939 \$4697 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10486 \$153 \$5070 \$5039 \$3731 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10487 \$153 \$5040 \$3651 \$5015 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10488 \$16 \$3852 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10489 \$153 \$4988 \$5041 \$3731 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10491 \$153 \$4988 \$3788 \$5016 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10492 \$16 \$3791 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10495 \$16 \$4949 \$4881 \$4989 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$10496 \$16 \$3792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10497 \$153 \$4950 \$4698 \$3792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10498 \$153 \$4990 \$5042 \$3852 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10499 \$153 \$4990 \$3763 \$4951 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10500 \$16 \$3731 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10501 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$10502 \$16 \$3852 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10504 \$153 \$5071 \$4931 \$3852 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10505 \$153 \$4991 \$3788 \$4992 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10506 \$153 \$5072 \$4952 \$3852 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10507 \$16 \$4882 \$4724 \$4932 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$10509 \$153 \$4910 \$3939 \$4639 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10511 \$153 \$4995 \$4920 \$3852 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10512 \$153 \$4995 \$3763 \$4953 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10513 \$16 \$4837 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10514 \$16 \$3731 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10515 \$16 \$4837 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10516 \$16 \$5158 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10517 \$16 \$3852 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10518 \$153 \$4998 \$5043 \$3852 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10520 \$16 \$5235 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10521 \$16 \$3852 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10523 \$153 \$5073 \$4804 \$3852 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10525 \$16 \$3731 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10527 \$16 \$3791 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10528 \$153 \$4804 \$4831 \$5000 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$10529 \$153 \$4955 \$4804 \$4048 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10530 \$16 \$4347 \$16 \$153 \$4937 VNB sky130_fd_sc_hd__clkbuf_2
X$10532 \$16 \$4317 \$16 \$153 \$5001 VNB sky130_fd_sc_hd__clkbuf_2
X$10533 \$16 \$5044 \$16 \$153 \$4834 VNB sky130_fd_sc_hd__clkbuf_2
X$10534 \$153 \$4956 \$4833 \$4935 \$4912 \$4933 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$10535 \$153 \$4912 \$4833 \$5018 \$4933 \$4935 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$10536 \$16 \$5018 \$16 \$153 \$5017 VNB sky130_fd_sc_hd__clkbuf_2
X$10538 \$16 \$5074 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10539 \$153 \$5045 \$4936 \$4958 \$5001 \$4937 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$10540 \$16 \$4834 \$16 \$153 \$4807 VNB sky130_fd_sc_hd__inv_1
X$10541 \$153 \$4964 \$3719 \$4963 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10543 \$153 \$5075 \$4887 \$3721 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10544 \$16 \$4921 \$16 \$153 \$4837 VNB sky130_fd_sc_hd__clkbuf_2
X$10545 \$16 \$3721 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10546 \$153 \$5004 \$4887 \$3691 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10547 \$153 \$4888 \$4414 \$4807 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10548 \$153 \$5093 \$3719 \$5019 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10550 \$153 \$4922 \$3986 \$4807 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10551 \$153 \$4960 \$3565 \$4807 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10552 \$153 \$4962 \$4626 \$3691 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10553 \$16 \$5017 \$16 \$153 \$4484 VNB sky130_fd_sc_hd__inv_1
X$10554 \$16 \$4949 \$5116 \$5020 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$10555 \$153 \$4627 \$4756 \$5020 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$10557 \$153 \$5005 \$3893 \$4484 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10559 \$153 \$5076 \$4627 \$3680 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10560 \$16 \$4949 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10561 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$10562 \$16 \$3898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10563 \$153 \$4890 \$4627 \$3898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10564 \$16 \$3680 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10565 \$16 \$4057 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10566 \$16 \$3602 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10568 \$16 \$4882 \$4736 \$5006 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$10569 \$16 \$3680 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10570 \$153 \$5003 \$4737 \$4057 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10571 \$16 \$3721 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10572 \$16 \$4882 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10573 \$16 \$3721 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10574 \$153 \$5265 \$4737 \$3721 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10575 \$153 \$4287 \$3719 \$4857 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10576 \$16 \$4803 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10578 \$153 \$4573 \$3142 \$4857 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10579 \$16 \$3691 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10581 \$153 \$4915 \$3676 \$4646 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10582 \$153 \$5008 \$3142 \$4646 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10583 \$16 \$3680 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10584 \$16 \$3680 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10585 \$16 \$4831 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10586 \$153 \$4740 \$4831 \$5009 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$10587 \$16 \$4830 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10589 \$16 \$3680 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10591 \$153 \$4964 \$4892 \$3680 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10592 \$16 \$3826 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10593 \$153 \$5046 \$3676 \$4965 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10594 \$153 \$5012 \$4892 \$3826 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10596 \$16 \$3898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10597 \$153 \$4521 \$3860 \$4537 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10599 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$10600 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$10601 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$10603 \$153 \$5077 \$4864 \$3616 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10604 \$153 \$5077 \$3389 \$4859 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10606 \$153 \$5104 \$5055 \$5120 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10607 \$16 \$4902 \$4538 \$5121 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$10608 \$153 \$5078 \$4864 \$3571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10609 \$153 \$5078 \$3422 \$4859 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10610 \$16 \$3571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10611 \$16 \$4742 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10613 \$153 \$5047 \$3422 \$4692 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10614 \$16 \$3571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10617 \$153 \$4788 \$5314 \$5049 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$10618 \$153 \$4614 \$5051 \$5050 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$10619 \$153 \$5079 \$4614 \$3616 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10620 \$153 \$5079 \$3389 \$4707 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10621 \$16 \$3616 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10624 \$16 \$5051 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10626 \$153 \$5052 \$3394 \$4693 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10627 \$153 \$5105 \$4789 \$3616 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10629 \$153 \$4971 \$3478 \$4693 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10630 \$16 \$3616 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10631 \$153 \$5081 \$4865 \$3571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10633 \$153 \$5081 \$3422 \$4940 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10634 \$16 \$4947 \$16 \$153 \$4940 VNB sky130_fd_sc_hd__inv_1
X$10635 \$153 \$5123 \$4865 \$3616 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10636 \$16 \$4947 \$4538 \$5122 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$10638 \$153 \$5024 \$4867 \$3571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10639 \$16 \$3571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10640 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$10642 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$10644 \$153 \$4709 \$4867 \$3616 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10645 \$16 \$5026 \$4012 \$5124 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$10646 \$153 \$5082 \$4791 \$3616 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10647 \$153 \$5082 \$3389 \$4941 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10648 \$16 \$3616 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10649 \$16 \$3571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10652 \$153 \$5056 \$3478 \$4941 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10653 \$153 \$5057 \$3394 \$4941 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10654 \$16 \$5184 \$5095 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$10655 \$153 \$5025 \$4711 \$3571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10656 \$16 \$5106 \$4631 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$10657 \$153 \$5126 \$4711 \$3616 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10659 \$16 \$3616 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10661 \$16 \$4706 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10662 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10663 \$153 \$3779 \$1482 \$5107 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10664 \$16 \$5107 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10666 \$16 \$5059 \$16 \$153 \$4822 VNB sky130_fd_sc_hd__clkbuf_2
X$10667 \$16 \$5058 \$16 \$153 \$3658 VNB sky130_fd_sc_hd__clkbuf_2
X$10668 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10669 \$16 \$5027 \$16 \$153 \$4893 VNB sky130_fd_sc_hd__clkbuf_2
X$10670 \$153 \$5128 \$4079 \$5127 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$10671 \$16 \$4275 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10673 \$16 \$4902 \$4275 \$5028 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$10674 \$16 \$6451 \$16 \$153 \$3241 VNB sky130_fd_sc_hd__clkbuf_2
X$10675 \$16 \$6451 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10677 \$153 \$5083 \$4926 \$3572 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10678 \$153 \$5083 \$3101 \$4861 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10679 \$16 \$3572 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10681 \$153 \$4750 \$3079 \$4529 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10682 \$16 \$5151 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10683 \$16 \$3692 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10685 \$16 \$5080 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10687 \$153 \$5030 \$4926 \$3492 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10688 \$153 \$4816 \$3354 \$4529 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10689 \$16 \$3492 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10690 \$153 \$5032 \$4873 \$3572 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10691 \$153 \$5108 \$3556 \$4796 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10692 \$16 \$3572 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10693 \$16 \$4939 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10695 \$153 \$4797 \$4939 \$5229 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$10696 \$16 \$3480 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10697 \$153 \$5035 \$4797 \$3480 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10698 \$16 \$3480 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10699 \$16 \$4893 \$4275 \$5129 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$10701 \$153 \$4927 \$4797 \$3543 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10704 \$16 \$3572 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10705 \$153 \$5062 \$3101 \$4818 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10707 \$16 \$4947 \$4275 \$5130 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$10708 \$153 \$5036 \$4622 \$3572 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10709 \$16 \$3572 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10710 \$16 \$4275 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10712 \$153 \$5014 \$4875 \$3543 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10715 \$153 \$5084 \$4875 \$3572 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10716 \$153 \$5084 \$3101 \$4798 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10718 \$153 \$4876 \$5109 \$5064 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$10719 \$153 \$5131 \$4876 \$3543 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10721 \$153 \$5038 \$4876 \$3572 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10722 \$16 \$4822 \$3957 \$5132 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$10723 \$16 \$3572 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10725 \$153 \$5085 \$4948 \$3572 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10726 \$153 \$5085 \$3101 \$5066 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10727 \$16 \$4983 \$16 \$153 \$3344 VNB sky130_fd_sc_hd__clkbuf_2
X$10729 \$16 \$3310 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10731 \$153 \$3310 \$3241 \$4620 \$3344 \$16 \$16 VNB sky130_fd_sc_hd__nor3b_4
X$10732 \$153 \$153 \$5096 \$5155 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10733 \$153 \$5067 \$3504 \$5066 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10735 \$153 \$4223 \$1482 \$5205 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10736 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10737 \$16 \$5096 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10738 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10740 \$153 \$3576 \$1482 \$5096 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10741 \$153 \$5133 \$4799 \$4048 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10742 \$153 \$5097 \$5110 \$3731 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10743 \$16 \$3791 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10744 \$16 \$3814 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10745 \$16 \$4760 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10746 \$16 \$3852 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10748 \$153 \$5134 \$5110 \$3852 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10749 \$16 \$3731 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10750 \$16 \$3852 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10751 \$153 \$5135 \$5039 \$3852 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10752 \$16 \$3731 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10753 \$153 \$5135 \$3763 \$5015 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10754 \$153 \$5111 \$3939 \$5015 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10756 \$153 \$5086 \$5041 \$3852 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10757 \$153 \$5086 \$3763 \$5016 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10758 \$16 \$3814 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10759 \$16 \$3791 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10760 \$153 \$5087 \$5042 \$3791 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10761 \$153 \$5087 \$3919 \$4951 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10762 \$16 \$3852 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10764 \$153 \$5088 \$5042 \$3731 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10765 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$10766 \$16 \$3791 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10767 \$153 \$5136 \$4931 \$3791 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10768 \$153 \$5071 \$3763 \$4992 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10770 \$153 \$4908 \$3939 \$4587 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10772 \$153 \$5137 \$4952 \$3791 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10773 \$153 \$5072 \$3763 \$5138 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10775 \$16 \$3852 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10777 \$153 \$5089 \$4920 \$3791 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10778 \$153 \$5089 \$3919 \$4953 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10779 \$16 \$3791 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10781 \$153 \$5090 \$5043 \$3791 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10783 \$16 \$3792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10784 \$16 \$3852 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10785 \$153 \$4998 \$3763 \$5139 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10787 \$153 \$5091 \$5112 \$3852 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10788 \$153 \$4999 \$3962 \$4700 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10790 \$153 \$5091 \$3763 \$5113 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10791 \$153 \$5092 \$5112 \$3791 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10792 \$153 \$5092 \$3919 \$5113 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10793 \$16 \$5355 \$5002 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$10794 \$153 \$5044 \$4933 \$4935 \$4912 \$4833 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$10795 \$153 \$4997 \$3676 \$4954 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10797 \$16 \$4935 \$4833 \$4912 \$4933 \$16 \$153 \$5140 VNB
+ sky130_fd_sc_hd__and4_2
X$10798 \$153 \$4936 \$5001 \$5141 \$4937 \$4958 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$10799 \$16 \$4930 \$5116 \$4886 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$10801 \$153 \$5098 \$3565 \$4963 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10802 \$153 \$5003 \$4414 \$3567 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10803 \$153 \$5075 \$3676 \$4807 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10804 \$16 \$5141 \$16 \$153 \$4830 VNB sky130_fd_sc_hd__clkbuf_2
X$10805 \$16 \$4057 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10807 \$153 \$5142 \$4414 \$5114 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10808 \$16 \$3691 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10809 \$153 \$5115 \$3565 \$5114 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10810 \$153 \$5093 \$5197 \$3680 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10812 \$16 \$5017 \$5116 \$5099 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$10813 \$153 \$4626 \$5498 \$5099 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$10816 \$16 \$3691 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10817 \$153 \$4913 \$3860 \$4484 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10818 \$153 \$5100 \$3565 \$5019 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10819 \$16 \$4756 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10820 \$16 \$5498 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10821 \$16 \$5017 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10822 \$153 \$5101 \$3719 \$5117 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10823 \$153 \$5143 \$3565 \$5117 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10824 \$16 \$3680 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10825 \$153 \$5118 \$4414 \$5117 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10827 \$153 \$5221 \$3676 \$5117 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10828 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$10829 \$153 \$5102 \$4414 \$5119 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10830 \$153 \$5094 \$5198 \$3680 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10831 \$153 \$5094 \$3719 \$5119 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10833 \$153 \$4353 \$4414 \$4857 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10835 \$153 \$4516 \$3565 \$4857 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10836 \$153 \$4885 \$5163 \$3680 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10837 \$153 \$4354 \$3860 \$4857 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10838 \$16 \$5353 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10839 \$16 \$5353 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10840 \$153 \$4838 \$3986 \$5011 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10841 \$153 \$4840 \$3893 \$5011 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10843 \$153 \$5145 \$5144 \$3680 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10844 \$153 \$4765 \$4414 \$4646 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10845 \$16 \$3691 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10846 \$16 \$3680 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10847 \$16 \$4057 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10848 \$153 \$5103 \$3719 \$4965 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10849 \$153 \$5146 \$4892 \$4057 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10851 \$16 \$3721 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10852 \$153 \$5147 \$4892 \$3721 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10853 \$153 \$7455 \$4892 \$3898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10854 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$10856 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$10857 \$153 \$950 \$234 \$783 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10858 \$153 \$967 \$816 \$263 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10859 \$153 \$921 \$102 \$763 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10860 \$153 \$968 \$816 \$58 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10861 \$16 \$58 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10864 \$16 \$945 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10865 \$153 \$969 \$816 \$184 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10866 \$153 \$869 \$349 \$763 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10867 \$16 \$184 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10868 \$16 \$419 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10869 \$153 \$951 \$349 \$1012 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10870 \$153 \$970 \$952 \$395 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10872 \$16 \$395 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10873 \$16 \$1291 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10874 \$16 \$1263 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10875 \$153 \$953 \$59 \$783 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10876 \$16 \$184 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10878 \$153 \$971 \$952 \$419 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10879 \$16 \$419 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10880 \$16 \$1013 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10881 \$16 \$972 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10882 \$153 \$954 \$755 \$263 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10885 \$153 \$714 \$102 \$903 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10887 \$16 \$419 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10888 \$153 \$973 \$817 \$249 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10889 \$153 \$954 \$234 \$903 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10890 \$153 \$924 \$102 \$639 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10891 \$153 \$973 \$377 \$639 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10893 \$153 \$840 \$394 \$639 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10894 \$153 \$871 \$234 \$765 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10895 \$153 \$974 \$664 \$504 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10896 \$16 \$504 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10897 \$16 \$1659 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10898 \$16 \$1594 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10899 \$153 \$975 \$756 \$395 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10902 \$153 \$841 \$59 \$651 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10904 \$153 \$976 \$756 \$263 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10905 \$153 \$873 \$349 \$651 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10906 \$153 \$976 \$234 \$651 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10907 \$16 \$652 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10908 \$153 \$874 \$234 \$766 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10911 \$153 \$977 \$1038 \$249 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10913 \$153 \$460 \$561 \$173 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10914 \$153 \$925 \$955 \$504 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10915 \$153 \$925 \$561 \$906 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10916 \$16 \$504 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10917 \$16 \$17 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10919 \$153 \$978 \$955 \$17 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10920 \$16 \$280 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10922 \$16 \$1037 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10923 \$16 \$979 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10924 \$153 \$820 \$819 \$187 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10926 \$16 \$1037 \$16 \$153 \$810 VNB sky130_fd_sc_hd__inv_1
X$10927 \$153 \$926 \$346 \$810 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10928 \$16 \$187 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10929 \$16 \$293 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10931 \$153 \$980 \$819 \$358 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10932 \$16 \$358 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10933 \$153 \$907 \$819 \$60 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10934 \$153 \$927 \$347 \$810 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10936 \$16 \$212 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10939 \$16 \$73 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10940 \$16 \$981 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10941 \$16 \$358 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10943 \$153 \$928 \$104 \$767 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10944 \$16 \$972 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10946 \$16 \$582 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10947 \$153 \$982 \$956 \$358 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10948 \$16 \$358 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10949 \$153 \$983 \$956 \$187 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10951 \$153 \$984 \$956 \$293 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10952 \$153 \$985 \$823 \$60 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10953 \$153 \$324 \$347 \$186 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10954 \$153 \$404 \$35 \$186 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10955 \$16 \$849 \$555 \$929 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$10958 \$153 \$986 \$900 \$18 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10959 \$16 \$209 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10961 \$153 \$987 \$900 \$73 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10962 \$153 \$988 \$900 \$358 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10963 \$16 \$899 \$507 \$930 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$10965 \$16 \$60 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10966 \$153 \$851 \$35 \$655 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10967 \$153 \$848 \$253 \$1040 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10968 \$16 \$293 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10969 \$16 \$1659 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10970 \$16 \$899 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10971 \$153 \$989 \$957 \$73 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10972 \$153 \$989 \$215 \$910 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10973 \$16 \$716 \$946 \$931 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$10975 \$153 \$990 \$957 \$60 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10976 \$16 \$209 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10977 \$153 \$991 \$759 \$73 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10978 \$153 \$991 \$215 \$760 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10979 \$153 \$932 \$35 \$760 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10980 \$16 \$209 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10981 \$16 \$18 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10983 \$153 \$933 \$253 \$760 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10984 \$153 \$852 \$389 \$656 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10985 \$16 \$424 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10987 \$16 \$902 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10989 \$16 \$145 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10990 \$16 \$1459 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$10991 \$153 \$826 \$1459 \$1015 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$10992 \$153 \$934 \$559 \$947 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10993 \$16 \$902 \$16 \$153 \$656 VNB sky130_fd_sc_hd__inv_1
X$10995 \$153 \$994 \$854 \$424 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$10996 \$153 \$935 \$559 \$656 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$10998 \$153 \$992 \$21 \$656 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11000 \$16 \$241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11001 \$153 \$995 \$590 \$241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11002 \$153 \$995 \$388 \$605 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11005 \$16 \$273 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11006 \$153 \$959 \$44 \$813 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11007 \$153 \$996 \$958 \$273 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11008 \$153 \$996 \$389 \$813 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11009 \$153 \$696 \$353 \$913 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11010 \$16 \$145 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11011 \$153 \$697 \$389 \$913 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11013 \$153 \$670 \$998 \$960 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$11014 \$153 \$997 \$559 \$814 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11015 \$153 \$961 \$266 \$814 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11016 \$153 \$1000 \$592 \$145 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11017 \$16 \$145 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11018 \$16 \$948 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11019 \$16 \$268 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11020 \$16 \$901 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11022 \$16 \$901 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11023 \$16 \$815 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11024 \$16 \$441 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11025 \$16 \$241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11026 \$153 \$962 \$21 \$1057 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11027 \$153 \$1001 \$1043 \$241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11028 \$153 \$1001 \$388 \$1057 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11029 \$153 \$999 \$21 \$1456 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11030 \$16 \$815 \$441 \$914 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$11032 \$153 \$938 \$893 \$424 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11033 \$16 \$724 \$441 \$894 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$11034 \$153 \$672 \$830 \$79 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11037 \$16 \$145 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11038 \$153 \$963 \$266 \$915 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11040 \$153 \$917 \$761 \$310 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11041 \$153 \$1002 \$761 \$446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11042 \$153 \$1002 \$393 \$774 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11045 \$153 \$939 \$761 \$309 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11046 \$16 \$309 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11047 \$16 \$309 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11048 \$153 \$896 \$596 \$509 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11049 \$16 \$964 \$16 \$153 \$658 VNB sky130_fd_sc_hd__inv_1
X$11050 \$153 \$1003 \$596 \$309 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11053 \$153 \$1003 \$703 \$658 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11054 \$16 \$446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11055 \$153 \$965 \$762 \$446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11057 \$16 \$63 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11058 \$153 \$1004 \$762 \$149 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11059 \$153 \$965 \$393 \$659 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11062 \$153 \$1005 \$706 \$446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11063 \$153 \$833 \$706 \$63 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11065 \$16 \$948 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11066 \$16 \$310 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11067 \$153 \$1007 \$1006 \$310 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11070 \$153 \$1007 \$223 \$949 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11073 \$153 \$1017 \$703 \$949 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11074 \$16 \$149 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11075 \$16 \$446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11076 \$153 \$751 \$943 \$149 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11078 \$16 \$309 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11079 \$153 \$865 \$371 \$779 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11080 \$153 \$918 \$966 \$509 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11082 \$153 \$1136 \$703 \$898 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11083 \$16 \$724 \$16 \$153 \$779 VNB sky130_fd_sc_hd__inv_1
X$11085 \$153 \$1010 \$966 \$178 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11086 \$16 \$178 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11087 \$153 \$1011 \$23 \$898 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11088 \$153 \$944 \$398 \$779 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11091 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$11092 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$11093 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$11094 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$11095 \$153 \$1045 \$234 \$1012 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11096 \$153 \$1018 \$394 \$1012 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11098 \$16 \$263 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11099 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$11100 \$153 \$1018 \$1036 \$395 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11101 \$153 \$968 \$30 \$763 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11102 \$16 \$395 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11104 \$16 \$249 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11105 \$153 \$816 \$945 \$1064 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$11106 \$16 \$1037 \$16 \$153 \$763 VNB sky130_fd_sc_hd__inv_1
X$11107 \$16 \$981 \$16 \$153 \$1012 VNB sky130_fd_sc_hd__inv_1
X$11110 \$153 \$1065 \$1036 \$184 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11111 \$16 \$184 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11112 \$153 \$953 \$952 \$184 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11113 \$153 \$950 \$952 \$263 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11114 \$16 \$263 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11115 \$16 \$58 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11116 \$16 \$1013 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11118 \$153 \$1046 \$377 \$783 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11119 \$153 \$971 \$349 \$783 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11120 \$153 \$1066 \$755 \$395 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11121 \$16 \$395 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11122 \$16 \$263 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11123 \$16 \$279 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11124 \$153 \$1019 \$817 \$184 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11126 \$16 \$184 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11128 \$153 \$1020 \$817 \$58 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11129 \$153 \$1020 \$30 \$639 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11130 \$16 \$899 \$537 \$1021 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$11131 \$153 \$664 \$1659 \$1021 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$11132 \$153 \$872 \$394 \$765 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11134 \$16 \$17 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11135 \$153 \$974 \$561 \$765 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11136 \$16 \$1067 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11137 \$16 \$899 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11138 \$153 \$756 \$1047 \$904 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$11139 \$16 \$395 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11140 \$16 \$1047 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11141 \$153 \$1022 \$1118 \$504 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11142 \$16 \$504 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11143 \$16 \$1264 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11145 \$16 \$1264 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11147 \$16 \$263 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11148 \$16 \$1048 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11149 \$153 \$1068 \$1038 \$419 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11150 \$16 \$419 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11152 \$16 \$504 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11153 \$153 \$1069 \$1038 \$504 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11154 \$16 \$249 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11155 \$16 \$1508 \$16 \$153 \$1070 VNB sky130_fd_sc_hd__inv_1
X$11157 \$153 \$284 \$234 \$173 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11159 \$153 \$905 \$955 \$263 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11160 \$16 \$419 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11161 \$16 \$263 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11163 \$16 \$395 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11164 \$153 \$1071 \$955 \$395 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11165 \$16 \$945 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11166 \$153 \$819 \$945 \$1072 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$11169 \$153 \$1073 \$1039 \$293 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11170 \$153 \$845 \$35 \$810 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11172 \$153 \$1074 \$1039 \$358 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11173 \$153 \$980 \$253 \$810 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11174 \$16 \$358 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11175 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$11177 \$16 \$212 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11179 \$16 \$1208 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11180 \$16 \$60 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11181 \$153 \$1075 \$758 \$212 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11182 \$153 \$1023 \$758 \$209 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11183 \$153 \$1023 \$346 \$767 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11184 \$16 \$209 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11185 \$16 \$1013 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11186 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$11188 \$153 \$1049 \$956 \$212 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11189 \$16 \$209 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11190 \$153 \$1076 \$956 \$73 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11191 \$16 \$73 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11193 \$153 \$290 \$54 \$186 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11194 \$153 \$403 \$253 \$186 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11197 \$153 \$1014 \$823 \$73 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11198 \$153 \$982 \$253 \$1111 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11199 \$16 \$73 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11200 \$153 \$1024 \$900 \$60 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11201 \$153 \$1024 \$104 \$909 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11202 \$16 \$60 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11203 \$16 \$293 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11206 \$153 \$987 \$215 \$909 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11207 \$153 \$1077 \$1041 \$60 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11208 \$153 \$1078 \$1041 \$73 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11209 \$16 \$73 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11211 \$16 \$18 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11213 \$153 \$891 \$957 \$18 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11214 \$16 \$73 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11216 \$153 \$1079 \$957 \$358 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11217 \$153 \$990 \$104 \$910 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11218 \$153 \$1079 \$253 \$910 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11219 \$16 \$60 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11222 \$16 \$1139 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11224 \$16 \$187 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11225 \$16 \$73 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11226 \$153 \$1050 \$54 \$1051 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11228 \$153 \$1080 \$1042 \$209 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11229 \$153 \$1025 \$1042 \$18 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11230 \$16 \$212 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11231 \$16 \$1551 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11232 \$16 \$241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11236 \$153 \$1081 \$1026 \$145 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11238 \$16 \$902 \$397 \$1015 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$11239 \$153 \$1082 \$1026 \$82 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11240 \$16 \$82 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11241 \$16 \$397 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11242 \$16 \$145 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11244 \$153 \$1027 \$854 \$145 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11245 \$153 \$1052 \$112 \$947 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11246 \$153 \$1083 \$854 \$82 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11247 \$153 \$855 \$388 \$657 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11249 \$16 \$964 \$397 \$1028 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$11251 \$153 \$590 \$884 \$1028 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$11252 \$16 \$82 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11253 \$153 \$959 \$958 \$82 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11254 \$153 \$1053 \$388 \$813 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11255 \$16 \$798 \$397 \$1054 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$11257 \$153 \$936 \$388 \$913 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11259 \$153 \$1055 \$112 \$813 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11261 \$16 \$901 \$268 \$960 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$11263 \$16 \$145 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11264 \$153 \$961 \$1056 \$145 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11265 \$16 \$273 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11267 \$153 \$1084 \$1056 \$273 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11268 \$16 \$829 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11269 \$16 \$998 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11270 \$16 \$82 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11271 \$153 \$1029 \$1043 \$82 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11272 \$153 \$1029 \$44 \$1057 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11273 \$153 \$1300 \$112 \$1412 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11275 \$153 \$1030 \$1043 \$145 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11276 \$153 \$1030 \$266 \$1057 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11278 \$153 \$1031 \$893 \$273 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11279 \$16 \$79 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11280 \$153 \$1031 \$389 \$915 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11281 \$16 \$79 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11284 \$153 \$1085 \$893 \$79 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11285 \$16 \$241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11286 \$153 \$1086 \$893 \$241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11287 \$153 \$963 \$893 \$145 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11288 \$16 \$902 \$369 \$1032 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$11291 \$153 \$761 \$1459 \$1032 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$11292 \$16 \$1044 \$16 \$153 \$1087 VNB sky130_fd_sc_hd__inv_1
X$11294 \$153 \$832 \$1058 \$149 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11295 \$16 \$964 \$369 \$1016 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$11298 \$153 \$1033 \$23 \$1087 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11300 \$153 \$550 \$371 \$258 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11302 \$153 \$1060 \$398 \$1059 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11303 \$153 \$762 \$998 \$940 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$11304 \$153 \$1061 \$23 \$1059 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11305 \$16 \$1062 \$16 \$153 \$369 VNB sky130_fd_sc_hd__clkbuf_2
X$11307 \$153 \$941 \$549 \$659 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11309 \$153 \$706 \$856 \$1034 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$11310 \$16 \$798 \$369 \$1034 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$11311 \$153 \$1063 \$223 \$1115 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11312 \$16 \$369 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11314 \$16 \$798 \$16 \$153 \$775 VNB sky130_fd_sc_hd__inv_1
X$11315 \$153 \$1005 \$393 \$775 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11316 \$16 \$856 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11320 \$16 \$149 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11321 \$16 \$446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11322 \$153 \$1035 \$1006 \$149 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11323 \$153 \$1035 \$398 \$949 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11325 \$153 \$1017 \$1006 \$309 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11327 \$153 \$1008 \$23 \$949 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11329 \$16 \$178 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11330 \$153 \$1088 \$943 \$178 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11331 \$16 \$509 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11332 \$153 \$1009 \$23 \$776 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11333 \$153 \$836 \$895 \$867 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$11336 \$153 \$1089 \$966 \$63 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11337 \$16 \$1120 \$16 \$153 \$898 VNB sky130_fd_sc_hd__inv_1
X$11338 \$16 \$509 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11340 \$16 \$149 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11341 \$153 \$919 \$966 \$149 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11342 \$153 \$1090 \$966 \$446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11344 \$153 \$920 \$966 \$310 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11345 \$16 \$310 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11346 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$11347 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$11348 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$11349 \$16 \$10427 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11350 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$11351 \$153 \$11732 \$10276 \$11717 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11352 \$153 \$11749 \$11733 \$10427 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11353 \$16 \$10295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11355 \$153 \$11750 \$11733 \$10646 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11356 \$16 \$10646 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11357 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$11360 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$11361 \$16 \$10427 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11362 \$153 \$11734 \$10705 \$11717 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11363 \$153 \$11683 \$11751 \$10427 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11364 \$153 \$11752 \$11751 \$10476 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11365 \$153 \$11683 \$10327 \$11718 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11368 \$153 \$11649 \$11631 \$10295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11369 \$16 \$10295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11370 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$11372 \$153 \$11753 \$11631 \$10368 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11373 \$153 \$11686 \$10327 \$11650 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11374 \$16 \$10368 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11375 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$11377 \$153 \$11754 \$11632 \$10476 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11378 \$16 \$10476 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11379 \$16 \$10427 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11380 \$153 \$11755 \$11632 \$10427 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11381 \$16 \$10427 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11382 \$153 \$11651 \$11633 \$10427 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11385 \$16 \$10368 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11386 \$16 \$10200 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11388 \$153 \$11756 \$11633 \$10476 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11389 \$16 \$10476 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11390 \$16 \$11897 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11392 \$16 \$10427 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11393 \$153 \$11687 \$11735 \$10427 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11394 \$153 \$11687 \$10327 \$11719 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11395 \$16 \$10476 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11398 \$153 \$11653 \$11735 \$10646 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11399 \$16 \$10646 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11401 \$16 \$10427 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11402 \$153 \$11688 \$11801 \$10427 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11403 \$153 \$11595 \$10276 \$11395 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11404 \$153 \$11688 \$10327 \$11655 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11406 \$153 \$11758 \$11801 \$10646 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11407 \$16 \$10368 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11408 \$16 \$10295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11410 \$153 \$11759 \$11429 \$11428 \$11430 \$11427 \$16 \$16 VNB
+ sky130_fd_sc_hd__nor4b_2
X$11411 \$16 \$11427 \$11430 \$11428 \$11429 \$16 \$153 \$11760 VNB
+ sky130_fd_sc_hd__and4_2
X$11412 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$11413 \$153 \$11736 \$11561 \$11529 \$11508 \$11507 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$11414 \$16 \$11720 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11416 \$153 \$11507 \$11561 \$11761 \$11508 \$11529 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$11417 \$16 \$11636 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11419 \$153 \$11656 \$11500 \$10606 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11420 \$153 \$11692 \$11737 \$10338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11421 \$153 \$11692 \$10309 \$11818 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11422 \$16 \$10338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11424 \$153 \$11762 \$11737 \$10470 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11425 \$16 \$10298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11426 \$16 \$10470 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11428 \$153 \$11763 \$11657 \$10338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11429 \$16 \$10338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11431 \$153 \$11693 \$11657 \$10298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11433 \$153 \$11763 \$10309 \$11838 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11434 \$16 \$10298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11435 \$16 \$11721 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11436 \$153 \$11764 \$11658 \$10338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11437 \$153 \$11659 \$11658 \$10298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11438 \$153 \$11764 \$10309 \$11562 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11439 \$16 \$10298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11441 \$153 \$11661 \$11967 \$10338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11442 \$16 \$11485 \$11164 \$11694 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$11443 \$16 \$10338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11444 \$153 \$11722 \$11967 \$10298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11445 \$153 \$11722 \$10401 \$11660 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11446 \$16 \$10298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11447 \$16 \$10382 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11448 \$16 \$11485 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11449 \$16 \$11897 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11451 \$16 \$11800 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11452 \$16 \$11800 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11453 \$16 \$10470 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11454 \$153 \$11738 \$10538 \$11488 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11455 \$153 \$11663 \$11639 \$10338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11456 \$153 \$11600 \$10344 \$11398 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11457 \$153 \$11664 \$11739 \$10298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11459 \$16 \$10298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11461 \$153 \$11765 \$11739 \$10338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11462 \$16 \$10338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11463 \$153 \$11575 \$11689 \$11740 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$11465 \$153 \$11576 \$11575 \$10298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11467 \$16 \$11594 \$16 \$153 \$11564 VNB sky130_fd_sc_hd__inv_1
X$11469 \$153 \$11766 \$10401 \$11488 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11470 \$153 \$11601 \$10098 \$11564 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11472 \$153 \$11767 \$11575 \$10605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11473 \$16 \$10338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11474 \$153 \$11697 \$10516 \$11564 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11475 \$153 \$11602 \$10247 \$11564 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11478 \$153 \$11768 \$11741 \$10300 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11479 \$16 \$10300 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11481 \$153 \$11769 \$11741 \$10611 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11482 \$153 \$11723 \$10919 \$11724 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11483 \$153 \$11770 \$10714 \$11724 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11485 \$16 \$10735 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11487 \$153 \$11771 \$11641 \$10735 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11488 \$16 \$10473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11489 \$16 \$11451 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11490 \$16 \$10809 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11491 \$153 \$11699 \$11666 \$10809 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11493 \$153 \$11699 \$10714 \$11513 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11495 \$16 \$11772 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11496 \$16 \$11772 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11497 \$16 \$10578 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11499 \$153 \$11579 \$11666 \$10578 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11500 \$153 \$11773 \$11742 \$10551 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11501 \$153 \$11643 \$11742 \$10473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11502 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$11504 \$16 \$11622 \$11378 \$11670 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$11505 \$153 \$11743 \$10919 \$11725 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11507 \$153 \$11744 \$10833 \$11725 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11508 \$153 \$11745 \$10471 \$11725 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11509 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$11511 \$16 \$10551 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11512 \$153 \$11774 \$11807 \$10551 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11514 \$16 \$10473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11515 \$16 \$10611 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11516 \$153 \$11775 \$11807 \$10611 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11517 \$16 \$11776 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11519 \$16 \$10551 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11520 \$153 \$11726 \$11645 \$10551 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11522 \$153 \$11726 \$10471 \$11727 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11524 \$16 \$11412 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11525 \$16 \$10735 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11527 \$153 \$11777 \$11645 \$10735 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11528 \$16 \$10611 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11529 \$16 \$10386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11530 \$153 \$11701 \$11580 \$10386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11531 \$16 \$10611 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11532 \$16 \$10735 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11533 \$153 \$11778 \$11580 \$10735 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11535 \$153 \$11779 \$11580 \$10809 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11536 \$153 \$11580 \$11747 \$11746 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$11537 \$16 \$11747 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11538 \$16 \$11459 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11539 \$16 \$11748 \$16 \$153 \$11502 VNB sky130_fd_sc_hd__clkbuf_2
X$11540 \$16 \$11147 \$16 \$153 \$11780 VNB sky130_fd_sc_hd__clkbuf_2
X$11541 \$16 \$11253 \$16 \$153 \$11781 VNB sky130_fd_sc_hd__clkbuf_2
X$11542 \$16 \$10986 \$16 \$153 \$11782 VNB sky130_fd_sc_hd__clkbuf_2
X$11543 \$16 \$11147 \$16 \$153 \$11582 VNB sky130_fd_sc_hd__clkbuf_2
X$11544 \$16 \$11374 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11546 \$16 \$11607 \$11646 \$11626 \$11582 \$16 \$153 \$11783 VNB
+ sky130_fd_sc_hd__and4_2
X$11547 \$153 \$11728 \$11582 \$11626 \$11646 \$11607 \$16 \$16 VNB
+ sky130_fd_sc_hd__nor4b_2
X$11548 \$153 \$11582 \$11646 \$11729 \$11626 \$11607 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$11549 \$16 \$11729 \$16 \$153 \$11172 VNB sky130_fd_sc_hd__clkbuf_2
X$11551 \$153 \$11784 \$11809 \$10326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11552 \$16 \$10326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11553 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$11555 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$11556 \$153 \$11704 \$11809 \$10393 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11557 \$153 \$11704 \$10694 \$11827 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11558 \$16 \$10393 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11559 \$153 \$11584 \$11628 \$10346 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11561 \$153 \$11705 \$10694 \$11829 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11563 \$16 \$10393 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11564 \$16 \$10346 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11566 \$153 \$11706 \$10694 \$11678 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11567 \$153 \$11785 \$11629 \$10564 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11569 \$16 \$11622 \$11504 \$11707 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$11570 \$153 \$11830 \$11629 \$10346 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11571 \$16 \$10346 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11572 \$16 \$10393 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11574 \$153 \$11679 \$11709 \$10326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11575 \$16 \$10326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11576 \$16 \$10446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11577 \$153 \$11786 \$11709 \$10446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11578 \$16 \$10326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11579 \$16 \$10346 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11580 \$153 \$11787 \$11681 \$10346 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11582 \$16 \$10446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11583 \$16 \$10393 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11584 \$153 \$11788 \$11681 \$10446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11585 \$153 \$11711 \$10694 \$11730 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11586 \$153 \$11788 \$10376 \$11730 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11587 \$16 \$10446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11588 \$153 \$11789 \$11587 \$10446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11590 \$16 \$10346 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11592 \$153 \$11712 \$10694 \$11731 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11593 \$16 \$11627 \$11229 \$11790 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$11595 \$153 \$11791 \$11588 \$10393 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11597 \$153 \$11868 \$11588 \$10326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11598 \$16 \$10393 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11599 \$16 \$11483 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11602 \$16 \$10326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11603 \$153 \$11387 \$10694 \$11461 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11604 \$153 \$11792 \$11648 \$10326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11606 \$16 \$10446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11607 \$153 \$11793 \$11648 \$10446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11608 \$153 \$11024 \$10376 \$11022 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11611 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$11612 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$11613 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$11614 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$11616 \$153 \$11732 \$11733 \$10295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11618 \$153 \$11749 \$10327 \$11717 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11620 \$153 \$11750 \$10318 \$11717 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11621 \$153 \$11734 \$11733 \$10476 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11622 \$16 \$10476 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11624 \$153 \$11811 \$11810 \$12150 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11625 \$153 \$11752 \$10705 \$11718 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11627 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$11629 \$153 \$11832 \$11751 \$10295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11631 \$153 \$11812 \$10330 \$11718 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11632 \$153 \$11684 \$10318 \$11718 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11634 \$153 \$11685 \$10705 \$11650 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11635 \$16 \$10226 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11636 \$16 \$10522 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11637 \$16 \$10539 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11639 \$16 \$10539 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11641 \$16 \$11794 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11642 \$16 \$10367 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11643 \$153 \$11753 \$10303 \$11650 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11644 \$16 \$11794 \$16 \$153 \$11650 VNB sky130_fd_sc_hd__inv_1
X$11645 \$16 \$11794 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11647 \$153 \$11568 \$11632 \$10295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11648 \$16 \$10295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11650 \$153 \$11754 \$10705 \$11560 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11651 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$11654 \$16 \$11721 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11655 \$153 \$11755 \$10327 \$11560 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11656 \$153 \$11615 \$11633 \$10200 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11658 \$153 \$11634 \$11633 \$10646 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11659 \$16 \$10646 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11660 \$153 \$11756 \$10705 \$11652 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11663 \$153 \$11833 \$11735 \$10476 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11664 \$153 \$11833 \$10705 \$11719 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11665 \$153 \$11992 \$10088 \$11719 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11666 \$16 \$10295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11667 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$11668 \$153 \$11813 \$10303 \$11719 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11669 \$16 \$10368 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11670 \$16 \$10367 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11671 \$16 \$11795 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11672 \$16 \$10476 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11674 \$153 \$11834 \$11801 \$10476 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11675 \$16 \$11814 \$16 \$153 \$11655 VNB sky130_fd_sc_hd__inv_1
X$11677 \$153 \$11654 \$11801 \$10295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11678 \$153 \$11758 \$10318 \$11655 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11679 \$16 \$11805 \$11689 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$11680 \$16 \$11815 \$16 \$153 \$11800 VNB sky130_fd_sc_hd__clkbuf_2
X$11681 \$16 \$11759 \$16 \$153 \$11795 VNB sky130_fd_sc_hd__clkbuf_2
X$11683 \$153 \$11815 \$11430 \$11427 \$11428 \$11429 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$11684 \$16 \$11529 \$11561 \$11508 \$11507 \$16 \$153 \$11835 VNB
+ sky130_fd_sc_hd__and4_2
X$11685 \$153 \$11508 \$11507 \$11816 \$11561 \$11529 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$11686 \$153 \$11508 \$11561 \$11836 \$11507 \$11529 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$11687 \$16 \$11636 \$11275 \$11691 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$11688 \$16 \$11761 \$16 \$153 \$11721 VNB sky130_fd_sc_hd__clkbuf_2
X$11689 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$11691 \$16 \$10606 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11693 \$16 \$10514 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11694 \$153 \$11817 \$10538 \$11818 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11695 \$153 \$11819 \$10686 \$11818 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11697 \$153 \$11837 \$11737 \$10298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11698 \$153 \$11837 \$10401 \$11818 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11699 \$153 \$11820 \$10098 \$11818 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11702 \$153 \$11762 \$10247 \$11818 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11703 \$16 \$11757 \$16 \$153 \$11838 VNB sky130_fd_sc_hd__inv_1
X$11705 \$153 \$11839 \$11657 \$10514 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11706 \$153 \$11839 \$10538 \$11838 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11707 \$153 \$11693 \$10401 \$11838 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11708 \$16 \$11757 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11709 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$11712 \$16 \$10338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11714 \$16 \$10514 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11715 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$11716 \$153 \$11840 \$11658 \$10382 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11717 \$153 \$11840 \$10098 \$11562 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11718 \$153 \$11662 \$11967 \$10470 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11719 \$16 \$10470 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11720 \$16 \$11164 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11722 \$16 \$10621 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11724 \$153 \$11638 \$11967 \$10382 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11725 \$16 \$10514 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11727 \$153 \$11204 \$11639 \$10470 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11728 \$16 \$11800 \$16 \$153 \$11488 VNB sky130_fd_sc_hd__inv_1
X$11730 \$153 \$11766 \$11639 \$10298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11733 \$16 \$10526 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11734 \$153 \$11821 \$10686 \$11563 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11735 \$153 \$11574 \$11739 \$10470 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11736 \$16 \$10526 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11737 \$16 \$10382 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11738 \$153 \$11640 \$11739 \$10382 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11739 \$153 \$11765 \$10309 \$11563 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11741 \$16 \$11594 \$11164 \$11740 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$11742 \$16 \$10298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11743 \$153 \$11841 \$11806 \$10298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11744 \$153 \$11695 \$10098 \$11488 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11745 \$16 \$10382 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11747 \$16 \$12476 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11748 \$16 \$10605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11749 \$153 \$11511 \$11806 \$10338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11752 \$153 \$11822 \$11806 \$10470 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11753 \$16 \$10470 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11754 \$153 \$11723 \$11741 \$10735 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11755 \$153 \$11796 \$11741 \$10473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11756 \$16 \$10473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11757 \$16 \$10386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11758 \$16 \$10809 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11760 \$153 \$11822 \$10247 \$11906 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11761 \$153 \$11823 \$10471 \$11724 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11762 \$153 \$11797 \$11641 \$10809 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11763 \$153 \$11796 \$10501 \$11724 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11764 \$153 \$11771 \$10919 \$11665 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11765 \$16 \$11824 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11766 \$16 \$10300 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11768 \$153 \$11490 \$11666 \$10300 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11769 \$16 \$11824 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11770 \$16 \$11842 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11771 \$16 \$10611 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11772 \$153 \$11843 \$11666 \$10611 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11773 \$16 \$10386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11774 \$153 \$11668 \$11742 \$10611 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11776 \$16 \$10809 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11777 \$16 \$10473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11778 \$153 \$11773 \$10471 \$11669 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11779 \$16 \$10473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11781 \$16 \$10735 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11782 \$153 \$11743 \$11880 \$10735 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11783 \$16 \$11622 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11785 \$16 \$10551 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11786 \$153 \$11745 \$11880 \$10551 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11788 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$11790 \$16 \$10735 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11791 \$153 \$11844 \$11807 \$10735 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11792 \$153 \$11845 \$11807 \$10473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11793 \$153 \$11774 \$10471 \$11954 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11794 \$16 \$11627 \$16 \$153 \$11954 VNB sky130_fd_sc_hd__inv_1
X$11796 \$16 \$10473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11797 \$16 \$10809 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11799 \$153 \$11671 \$11645 \$10473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11800 \$153 \$12049 \$10472 \$11727 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11802 \$16 \$11412 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11803 \$16 \$11798 \$16 \$153 \$11727 VNB sky130_fd_sc_hd__inv_1
X$11804 \$153 \$11777 \$10919 \$11727 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11805 \$153 \$11802 \$11808 \$10611 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11807 \$153 \$11674 \$11580 \$10611 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11808 \$153 \$11802 \$10833 \$11825 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11810 \$16 \$10300 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11811 \$153 \$11778 \$10919 \$11673 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11812 \$16 \$11412 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11813 \$16 \$11459 \$11412 \$11746 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$11814 \$153 \$11779 \$10714 \$11673 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11815 \$16 \$11459 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11818 \$16 \$11385 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11820 \$16 \$11826 \$16 \$153 \$11622 VNB sky130_fd_sc_hd__clkbuf_2
X$11821 \$153 \$11826 \$11780 \$11781 \$11782 \$11803 \$16 \$16 VNB
+ sky130_fd_sc_hd__nor4b_2
X$11822 \$16 \$11803 \$11782 \$11781 \$11780 \$16 \$153 \$11846 VNB
+ sky130_fd_sc_hd__and4_2
X$11824 \$16 \$11503 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11825 \$153 \$11847 \$11646 \$11607 \$11626 \$11582 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$11826 \$153 \$11626 \$11582 \$11848 \$11646 \$11607 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$11827 \$16 \$11728 \$16 \$153 \$11483 VNB sky130_fd_sc_hd__clkbuf_2
X$11828 \$16 \$11374 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11831 \$16 \$10564 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11832 \$153 \$11609 \$10815 \$11515 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11833 \$153 \$11702 \$10587 \$11515 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11834 \$153 \$11784 \$10466 \$11827 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11836 \$153 \$11849 \$11809 \$10346 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11837 \$153 \$11849 \$10285 \$11827 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11840 \$153 \$11828 \$10376 \$11827 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11841 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$11842 \$16 \$11016 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11844 \$153 \$11799 \$11628 \$10446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11845 \$153 \$11799 \$10376 \$11829 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11846 \$16 \$10564 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11847 \$16 \$10446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11849 \$153 \$11785 \$10642 \$11678 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11851 \$16 \$11622 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11853 \$16 \$10326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11854 \$153 \$11677 \$11629 \$10326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11855 \$153 \$11830 \$10285 \$11678 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11856 \$153 \$11850 \$10587 \$11678 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11857 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$11858 \$153 \$11708 \$10694 \$11680 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11859 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$11861 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$11862 \$16 \$10392 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11863 \$153 \$11710 \$10285 \$11680 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11864 \$153 \$11786 \$10376 \$11680 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11865 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$11866 \$153 \$11787 \$10285 \$11730 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11867 \$16 \$11413 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11868 \$16 \$12404 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11869 \$153 \$11587 \$12404 \$11804 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$11871 \$16 \$10467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11873 \$16 \$11413 \$11229 \$11804 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$11875 \$16 \$10617 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11876 \$153 \$11611 \$10466 \$11731 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11877 \$153 \$11851 \$11587 \$10617 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11878 \$153 \$11789 \$10376 \$11731 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11879 \$153 \$11831 \$10815 \$11731 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11880 \$16 \$10393 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11882 \$16 \$10326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11884 \$153 \$11517 \$10642 \$11390 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11885 \$16 \$10617 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11887 \$153 \$11852 \$11588 \$10467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11888 \$16 \$10467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11889 \$16 \$11390 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11891 \$16 \$11390 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11893 \$153 \$11324 \$10466 \$11461 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11894 \$153 \$10451 \$10466 \$10801 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11895 \$16 \$10446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11898 \$153 \$11853 \$11648 \$10467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11899 \$16 \$10467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11900 \$153 \$11110 \$10587 \$11022 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11901 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$11902 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$11903 \$153 \$12315 \$12412 \$12150 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11904 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$11905 \$153 \$12436 \$12229 \$12150 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11906 \$153 \$12467 \$12355 \$12152 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11907 \$153 \$12467 \$12209 \$12386 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11908 \$153 \$12437 \$12412 \$12386 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11909 \$16 \$12152 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11912 \$16 \$10764 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11913 \$16 \$12158 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11914 \$153 \$12250 \$12134 \$12020 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11916 \$153 \$12376 \$12355 \$12003 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11918 \$153 \$12438 \$12353 \$12386 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11919 \$153 \$12439 \$12229 \$12386 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11920 \$16 \$12095 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11921 \$16 \$10730 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11924 \$153 \$12468 \$12469 \$12003 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11925 \$16 \$12003 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11926 \$16 \$12158 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11927 \$153 \$12318 \$12412 \$12252 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11928 \$153 \$12469 \$11114 \$12387 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$11929 \$153 \$12793 \$12412 \$12563 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11930 \$16 \$11114 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11933 \$153 \$12440 \$12134 \$12426 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11934 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$11935 \$153 \$12441 \$11810 \$12426 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11937 \$153 \$12470 \$12471 \$12003 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11938 \$16 \$12003 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11940 \$153 \$12389 \$12412 \$12004 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11941 \$16 \$12095 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11942 \$16 \$8361 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11944 \$153 \$12471 \$11194 \$12442 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$11945 \$16 \$11194 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11947 \$153 \$12444 \$11993 \$12443 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$11948 \$16 \$12236 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11950 \$153 \$12472 \$12444 \$12093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11952 \$16 \$12003 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11953 \$16 \$10825 \$16 \$153 \$12413 VNB sky130_fd_sc_hd__inv_1
X$11955 \$153 \$12445 \$11810 \$12413 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11956 \$153 \$12390 \$12412 \$12005 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11957 \$153 \$12099 \$12172 \$12236 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11958 \$16 \$12236 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11959 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$11960 \$153 \$12414 \$12391 \$12003 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11962 \$16 \$12003 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11963 \$16 \$12095 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11964 \$153 \$12414 \$11810 \$12392 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11965 \$153 \$12473 \$12391 \$12093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11966 \$16 \$12294 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11967 \$16 \$12093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11969 \$16 \$10764 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11970 \$153 \$153 \$12209 \$12415 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11972 \$153 \$153 \$12353 \$12415 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11974 \$153 \$153 \$12134 \$12415 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11976 \$16 \$12295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11977 \$153 \$12416 \$12357 \$12296 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11978 \$153 \$12416 \$12359 \$12427 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11979 \$16 \$10764 \$16 \$153 \$12427 VNB sky130_fd_sc_hd__inv_1
X$11980 \$153 \$12417 \$12357 \$12101 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11982 \$153 \$12474 \$12357 \$12241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11983 \$153 \$12417 \$12476 \$12427 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11984 \$16 \$12241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11985 \$16 \$12241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11986 \$153 \$12475 \$12533 \$12083 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11987 \$153 \$12394 \$12363 \$12238 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11988 \$16 \$12083 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11990 \$153 \$12477 \$11114 \$12395 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$11992 \$153 \$12214 \$12363 \$12104 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11993 \$153 \$12478 \$12477 \$12295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$11994 \$153 \$12447 \$12028 \$12498 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$11995 \$16 \$12295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11997 \$16 \$12295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$11998 \$16 \$10722 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12000 \$153 \$12478 \$12155 \$12498 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12001 \$16 \$10825 \$12161 \$12479 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$12002 \$16 \$10825 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12004 \$153 \$12323 \$12359 \$12071 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12005 \$153 \$12396 \$12155 \$12071 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12006 \$153 \$12538 \$12028 \$12360 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12007 \$153 \$12448 \$12155 \$12360 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12008 \$16 \$11194 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12011 \$153 \$12480 \$12476 \$12360 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12012 \$153 \$12397 \$12363 \$12007 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12013 \$16 \$12296 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12014 \$153 \$11968 \$10344 \$11488 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12016 \$153 \$12428 \$12028 \$12429 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12017 \$16 \$12160 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12018 \$16 \$10624 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12019 \$16 \$11488 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12021 \$153 \$12398 \$12155 \$11869 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12024 \$153 \$12449 \$12359 \$12430 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12025 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$12026 \$153 \$12261 \$12363 \$11869 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12027 \$153 \$12450 \$12476 \$12430 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12029 \$153 \$12418 \$12308 \$12101 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12030 \$16 \$12101 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12031 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$12033 \$153 \$12418 \$12476 \$12378 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12034 \$16 \$16 \$153 VNB sky130_fd_sc_hd__conb_1
X$12035 \$16 \$10500 \$16 \$153 \$12431 VNB sky130_fd_sc_hd__clkbuf_2
X$12036 \$153 \$153 \$12476 \$12431 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12038 \$153 \$153 \$12174 \$12431 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12039 \$153 \$153 \$12155 \$12431 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12040 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$12042 \$16 \$12164 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12044 \$153 \$12419 \$12400 \$12164 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12045 \$153 \$12419 \$12217 \$12325 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12047 \$153 \$12420 \$12400 \$12298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12048 \$153 \$12420 \$12165 \$12325 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12049 \$16 \$12298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12051 \$16 \$12298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12053 \$153 \$12481 \$12482 \$12298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12054 \$16 \$11207 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12056 \$153 \$12482 \$11015 \$12401 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$12057 \$16 \$11015 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12058 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$12060 \$153 \$12328 \$12165 \$12216 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12061 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$12062 \$16 \$10739 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12063 \$16 \$10897 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12065 \$153 \$12402 \$12309 \$12216 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12067 \$153 \$12518 \$12347 \$12403 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$12068 \$153 \$12483 \$12309 \$12503 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12069 \$16 \$12347 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12070 \$16 \$11013 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12072 \$16 \$12571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12073 \$153 \$12310 \$12163 \$12571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12075 \$153 \$12421 \$12452 \$12326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12076 \$153 \$12453 \$12217 \$12432 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12077 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$12078 \$153 \$12454 \$12309 \$12432 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12079 \$16 \$12571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12080 \$153 \$12484 \$12113 \$12571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12083 \$153 \$12346 \$12217 \$12200 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12085 \$16 \$12164 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12086 \$16 \$12326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12087 \$153 \$12422 \$12075 \$12326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12088 \$153 \$12455 \$12603 \$11999 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12089 \$153 \$12422 \$12264 \$11999 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12091 \$16 \$12233 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12093 \$16 \$12571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12095 \$153 \$12485 \$12177 \$12571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12096 \$153 \$12456 \$12264 \$12117 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12098 \$16 \$12219 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12099 \$153 \$12486 \$12204 \$12219 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12101 \$153 \$12265 \$12165 \$12246 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12104 \$153 \$12487 \$12204 \$12164 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12105 \$16 \$12233 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12106 \$153 \$12381 \$12204 \$12233 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12108 \$16 \$12348 \$12404 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$12109 \$16 \$12348 \$11946 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$12110 \$16 \$10409 \$16 \$153 \$12488 VNB sky130_fd_sc_hd__inv_1
X$12111 \$16 \$10960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12112 \$16 \$12433 \$12009 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$12113 \$16 \$12168 \$16 \$153 \$12433 VNB sky130_fd_sc_hd__clkbuf_2
X$12114 \$16 \$12433 \$12198 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$12116 \$16 \$12433 \$12169 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$12117 \$16 \$11015 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12118 \$153 \$153 \$12339 \$12405 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12119 \$153 \$153 \$11942 \$12405 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12120 \$16 \$12348 \$11585 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$12121 \$153 \$12434 \$11015 \$12407 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$12122 \$16 \$12303 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12123 \$16 \$10978 \$16 \$153 \$12423 VNB sky130_fd_sc_hd__inv_1
X$12124 \$16 \$12299 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12125 \$153 \$12458 \$12119 \$12423 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12127 \$153 \$12382 \$12434 \$12303 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12128 \$153 \$12424 \$12434 \$12287 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12129 \$16 \$12287 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12131 \$16 \$11013 \$12459 \$12460 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$12132 \$153 \$12489 \$12347 \$12460 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$12133 \$16 \$12303 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12135 \$153 \$12424 \$12339 \$12423 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12136 \$16 \$12010 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12137 \$153 \$12461 \$12179 \$12337 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12139 \$153 \$12462 \$11942 \$12337 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12140 \$153 \$12463 \$12182 \$12337 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12141 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$12142 \$16 \$11622 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12143 \$153 \$12464 \$12339 \$12435 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12145 \$153 \$12465 \$12182 \$12435 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12147 \$16 \$12384 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12148 \$16 \$10552 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12149 \$153 \$12466 \$11942 \$12435 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12151 \$16 \$12299 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12152 \$153 \$12425 \$12180 \$12299 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12153 \$153 \$12425 \$12371 \$12302 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12154 \$16 \$12384 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12155 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$12157 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$12158 \$153 \$12268 \$11881 \$12302 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12160 \$16 \$12303 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12161 \$153 \$12408 \$12088 \$12303 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12162 \$153 \$12490 \$12088 \$12287 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12163 \$16 \$12245 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12164 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$12165 \$16 \$12303 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12167 \$153 \$12491 \$12409 \$12303 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12168 \$153 \$12492 \$12409 \$12351 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12169 \$16 \$10409 \$12018 \$12410 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$12171 \$153 \$12493 \$12373 \$11983 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12172 \$16 \$11983 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12174 \$16 \$10409 \$16 \$153 \$12411 VNB sky130_fd_sc_hd__inv_1
X$12175 \$153 \$12352 \$11942 \$12411 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12176 \$16 \$10409 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12178 \$16 \$12303 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12179 \$153 \$12385 \$12373 \$12303 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12180 \$153 \$12494 \$12373 \$12384 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12181 \$16 \$12384 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12182 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$12184 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$12185 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$12186 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$12187 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$12189 \$153 \$12437 \$12355 \$12230 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12191 \$16 \$12230 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12192 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$12193 \$153 \$12511 \$12208 \$12386 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12194 \$153 \$12522 \$12355 \$12158 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12195 \$153 \$12522 \$12057 \$12386 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12196 \$153 \$12439 \$12355 \$12093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12198 \$16 \$12093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12199 \$16 \$12003 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12200 \$16 \$11078 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12201 \$153 \$12513 \$11810 \$12512 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12202 \$16 \$10764 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12204 \$153 \$12523 \$12469 \$12093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12205 \$16 \$12093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12207 \$153 \$12524 \$12469 \$12158 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12210 \$16 \$10453 \$12012 \$12525 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$12211 \$153 \$12526 \$12586 \$12095 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12212 \$16 \$12095 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12213 \$16 \$10453 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12215 \$153 \$12527 \$12586 \$12093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12216 \$153 \$12527 \$12229 \$12426 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12217 \$16 \$12093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12218 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$12220 \$153 \$12528 \$12471 \$12095 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12221 \$153 \$12254 \$12134 \$12004 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12222 \$16 \$11077 \$12015 \$12442 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$12223 \$16 \$11077 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12224 \$153 \$12529 \$12471 \$12158 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12225 \$16 \$10825 \$12015 \$12443 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$12226 \$16 \$12158 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12229 \$16 \$10825 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12230 \$16 \$11993 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12232 \$153 \$12445 \$12444 \$12003 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12233 \$153 \$12472 \$12229 \$12413 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12235 \$16 \$10747 \$12015 \$12530 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$12236 \$153 \$12495 \$12514 \$12095 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12237 \$16 \$12095 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12240 \$153 \$12496 \$12514 \$12093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12241 \$16 \$10747 \$16 \$153 \$12579 VNB sky130_fd_sc_hd__inv_1
X$12242 \$16 \$12093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12243 \$16 \$10747 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12245 \$153 \$12531 \$12391 \$12095 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12246 \$153 \$12532 \$12391 \$12294 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12249 \$153 \$153 \$11810 \$12415 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12250 \$153 \$153 \$12057 \$12415 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12251 \$16 \$10500 \$16 \$153 \$12415 VNB sky130_fd_sc_hd__clkbuf_2
X$12252 \$153 \$12533 \$10634 \$12320 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$12254 \$16 \$12044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12255 \$153 \$12534 \$12357 \$12044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12257 \$153 \$12534 \$12068 \$12427 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12258 \$16 \$12259 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12259 \$16 \$12296 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12260 \$153 \$12497 \$12357 \$12160 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12261 \$153 \$12515 \$12174 \$12427 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12262 \$153 \$12497 \$12028 \$12427 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12263 \$153 \$12474 \$12363 \$12427 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12265 \$153 \$12535 \$12533 \$12160 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12266 \$153 \$12475 \$12174 \$12154 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12267 \$16 \$12160 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12268 \$16 \$10453 \$12159 \$12536 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$12269 \$153 \$12499 \$12477 \$12101 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12270 \$16 \$10939 \$16 \$153 \$12498 VNB sky130_fd_sc_hd__inv_1
X$12271 \$16 \$12101 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12272 \$16 \$10453 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12275 \$153 \$12537 \$12477 \$12083 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12276 \$16 \$12083 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12277 \$16 \$10939 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12279 \$16 \$11993 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12280 \$153 \$12500 \$11993 \$12479 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$12281 \$153 \$12538 \$12500 \$12160 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12282 \$16 \$12160 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12284 \$16 \$11077 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12285 \$16 \$11077 \$12161 \$12501 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$12286 \$153 \$12539 \$12500 \$12083 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12287 \$16 \$12083 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12289 \$153 \$12508 \$11194 \$12501 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$12290 \$153 \$12428 \$12508 \$12160 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12292 \$153 \$12502 \$10624 \$12509 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$12293 \$16 \$10747 \$12161 \$12509 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$12294 \$16 \$10747 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12295 \$16 \$10747 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12296 \$16 \$10747 \$16 \$153 \$12430 VNB sky130_fd_sc_hd__inv_1
X$12297 \$153 \$12540 \$12308 \$12295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12299 \$153 \$12540 \$12155 \$12378 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12300 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$12302 \$153 \$12541 \$12359 \$12378 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12303 \$153 \$12542 \$12308 \$12259 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12304 \$153 \$12542 \$12307 \$12378 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12305 \$16 \$12259 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12306 \$16 \$10500 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12307 \$153 \$153 \$12028 \$12431 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12308 \$153 \$153 \$12359 \$12431 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12310 \$153 \$153 \$12307 \$12431 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12311 \$153 \$153 \$12068 \$12431 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12313 \$16 \$12571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12314 \$16 \$12326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12315 \$153 \$12543 \$12400 \$12326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12317 \$153 \$12543 \$12264 \$12325 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12318 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$12321 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$12322 \$16 \$11113 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12323 \$16 \$11113 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12324 \$153 \$12516 \$12603 \$12325 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12326 \$16 \$12603 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12327 \$16 \$12264 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12328 \$16 \$12219 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12329 \$153 \$12544 \$12482 \$12219 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12330 \$153 \$12544 \$12110 \$12517 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12332 \$16 \$10978 \$16 \$153 \$12517 VNB sky130_fd_sc_hd__inv_1
X$12333 \$16 \$10978 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12336 \$16 \$12571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12337 \$16 \$12164 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12338 \$16 \$12115 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12339 \$153 \$12545 \$12482 \$12115 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12340 \$153 \$12545 \$12234 \$12517 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12342 \$153 \$12546 \$12518 \$12326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12343 \$16 \$12326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12345 \$16 \$12115 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12346 \$16 \$11013 \$16 \$153 \$12503 VNB sky130_fd_sc_hd__inv_1
X$12348 \$153 \$12547 \$12518 \$12115 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12349 \$16 \$10739 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12350 \$16 \$12115 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12351 \$16 \$12298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12352 \$16 \$12326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12353 \$153 \$12548 \$12452 \$12115 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12355 \$153 \$12548 \$12234 \$12432 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12356 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$12358 \$153 \$12421 \$12264 \$12432 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12359 \$16 \$12297 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12360 \$153 \$12549 \$12113 \$12297 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12361 \$153 \$12549 \$12582 \$12200 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12362 \$16 \$10552 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12363 \$16 \$12298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12364 \$153 \$12504 \$12075 \$12298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12366 \$153 \$12550 \$12075 \$12571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12367 \$16 \$12571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12368 \$16 \$12297 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12369 \$153 \$12551 \$12177 \$12297 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12370 \$153 \$12505 \$12177 \$12298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12371 \$16 \$12298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12372 \$16 \$12571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12374 \$153 \$12510 \$12204 \$12571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12376 \$153 \$12486 \$12110 \$12333 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12377 \$153 \$12510 \$12309 \$12333 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12378 \$16 \$10409 \$12166 \$12552 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$12379 \$153 \$12487 \$12217 \$12333 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12381 \$16 \$12348 \$11280 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$12382 \$16 \$12348 \$11921 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$12385 \$153 \$12519 \$12234 \$12333 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12386 \$153 \$12520 \$12264 \$12333 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12387 \$16 \$12326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12388 \$16 \$12433 \$11604 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$12389 \$16 \$10854 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12390 \$153 \$153 \$12119 \$12405 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12391 \$153 \$153 \$12371 \$12405 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12392 \$16 \$12348 \$11385 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$12393 \$153 \$153 \$12179 \$12405 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12396 \$153 \$12458 \$12434 \$12351 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12397 \$153 \$12553 \$12434 \$12299 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12398 \$16 \$12303 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12399 \$16 \$11113 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12401 \$16 \$12010 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12402 \$153 \$12554 \$12434 \$12010 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12404 \$16 \$12120 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12406 \$153 \$12288 \$12119 \$12247 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12407 \$153 \$12554 \$11942 \$12423 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12408 \$16 \$12384 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12409 \$153 \$12461 \$12489 \$12384 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12410 \$153 \$12462 \$12489 \$12010 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12413 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$12414 \$16 \$12287 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12415 \$16 \$12120 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12416 \$153 \$12465 \$12583 \$12120 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12417 \$16 \$11622 \$16 \$153 \$12435 VNB sky130_fd_sc_hd__inv_1
X$12418 \$153 \$12506 \$12583 \$12384 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12419 \$153 \$12506 \$12179 \$12435 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12420 \$16 \$10552 \$12018 \$12555 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$12422 \$153 \$12556 \$12180 \$12351 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12424 \$153 \$12557 \$12180 \$12384 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12425 \$153 \$12507 \$12180 \$12287 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12426 \$16 \$12287 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12427 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$12428 \$16 \$11413 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12430 \$153 \$12507 \$12339 \$12302 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12431 \$16 \$11983 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12433 \$16 \$12384 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12434 \$153 \$12558 \$12409 \$12384 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12435 \$16 \$11546 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12436 \$16 \$12010 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12437 \$153 \$12491 \$12227 \$12521 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12438 \$153 \$12558 \$12179 \$12521 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12439 \$16 \$12351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12440 \$16 \$10409 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12442 \$153 \$12492 \$12119 \$12521 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12443 \$16 \$12120 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12444 \$153 \$12559 \$12373 \$12120 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12445 \$153 \$12559 \$12182 \$12411 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12447 \$16 \$12299 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12448 \$153 \$12560 \$12373 \$12299 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12452 \$153 \$12560 \$12371 \$12411 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12453 \$153 \$12494 \$12179 \$12411 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12454 \$153 \$11853 \$10587 \$11926 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12455 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$12456 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$12457 \$153 \$7648 \$7544 \$6783 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12458 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$12459 \$16 \$6783 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12460 \$153 \$7649 \$7544 \$6784 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12461 \$153 \$7649 \$6794 \$7552 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12462 \$153 \$7618 \$6913 \$7552 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12463 \$16 \$6784 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12465 \$153 \$7650 \$7544 \$6792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12466 \$16 \$6792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12467 \$153 \$7544 \$7237 \$7619 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$12468 \$16 \$7545 \$7233 \$7619 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$12469 \$16 \$7237 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12470 \$153 \$7585 \$7053 \$6907 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12473 \$153 \$7585 \$6913 \$7137 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12474 \$16 \$6907 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12475 \$16 \$7521 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12476 \$153 \$7586 \$7620 \$6907 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12477 \$153 \$7586 \$6913 \$7587 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12478 \$16 \$6907 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12479 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$12481 \$153 \$7282 \$6719 \$7140 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12482 \$16 \$6981 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12484 \$153 \$7621 \$7546 \$6783 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12485 \$16 \$6783 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12487 \$153 \$7652 \$7546 \$6792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12488 \$16 \$6792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12490 \$153 \$7653 \$7546 \$7041 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12491 \$16 \$7041 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12493 \$153 \$7040 \$6930 \$6733 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12494 \$153 \$7653 \$6996 \$7608 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12495 \$153 \$7652 \$6719 \$7608 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12496 \$153 \$7588 \$7235 \$6792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12497 \$153 \$7588 \$6719 \$7142 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12498 \$16 \$6792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12499 \$16 \$6981 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12501 \$153 \$7651 \$6732 \$7609 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12502 \$16 \$6792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12503 \$16 \$6783 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12504 \$153 \$7654 \$7236 \$6783 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12506 \$153 \$7589 \$7337 \$6979 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12507 \$153 \$7589 \$6995 \$7439 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12510 \$16 \$6753 \$16 \$153 \$7439 VNB sky130_fd_sc_hd__inv_1
X$12511 \$153 \$7622 \$6913 \$7439 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12512 \$153 \$7286 \$6732 \$7437 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12513 \$16 \$7655 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12514 \$16 \$7590 \$16 \$153 \$7000 VNB sky130_fd_sc_hd__clkbuf_2
X$12515 \$153 \$7558 \$7472 \$7440 \$7456 \$7470 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$12516 \$153 \$7590 \$7470 \$7440 \$7456 \$7472 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$12517 \$16 \$7623 \$16 \$153 \$7072 VNB sky130_fd_sc_hd__clkbuf_2
X$12518 \$16 \$7381 \$6990 \$7591 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$12520 \$16 \$3384 \$16 \$153 \$7801 VNB sky130_fd_sc_hd__clkbuf_2
X$12521 \$16 \$4360 \$16 \$153 \$7656 VNB sky130_fd_sc_hd__clkbuf_2
X$12522 \$153 \$7657 \$7624 \$6862 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12523 \$153 \$7610 \$6992 \$7611 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12524 \$16 \$6862 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12525 \$16 \$7922 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12527 \$153 \$7404 \$7357 \$7044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12528 \$16 \$7060 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12530 \$153 \$7625 \$6756 \$7611 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12531 \$16 \$7044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12532 \$153 \$7626 \$6867 \$7611 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12533 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$12534 \$153 \$7658 \$7627 \$6991 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12536 \$153 \$7628 \$6324 \$7562 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12537 \$16 \$6991 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12538 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$12539 \$16 \$7521 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12542 \$16 \$7659 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12543 \$153 \$7629 \$6756 \$7562 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12544 \$16 \$7521 \$6990 \$7592 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$12546 \$16 \$7521 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12547 \$153 \$7660 \$7323 \$6771 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12548 \$16 \$6771 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12549 \$153 \$7661 \$7323 \$7060 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12550 \$16 \$6991 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12553 \$16 \$6916 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12554 \$153 \$7476 \$7335 \$7630 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$12555 \$153 \$7593 \$7476 \$6754 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12557 \$153 \$7593 \$6756 \$7458 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12558 \$153 \$7566 \$6867 \$7458 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12559 \$16 \$6754 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12560 \$16 \$7060 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12562 \$153 \$7685 \$7476 \$6771 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12563 \$153 \$7478 \$7238 \$6862 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12564 \$16 \$6862 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12565 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$12566 \$153 \$7662 \$7479 \$6916 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12567 \$16 \$6916 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12569 \$16 \$7663 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12570 \$16 \$6903 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12571 \$153 \$7594 \$7479 \$6991 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12572 \$153 \$7567 \$6906 \$7612 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12573 \$153 \$7594 \$6992 \$7612 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12574 \$153 \$7664 \$7006 \$7612 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12575 \$153 \$7568 \$6867 \$7411 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12577 \$16 \$6916 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12578 \$153 \$7569 \$6324 \$7411 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12579 \$153 \$7595 \$7708 \$7044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12581 \$153 \$7570 \$7003 \$7411 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12582 \$16 \$7044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12584 \$153 \$7256 \$7549 \$7082 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12586 \$153 \$7595 \$7006 \$7749 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12587 \$16 \$7386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12588 \$153 \$7631 \$7366 \$7296 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12589 \$153 \$7013 \$7347 \$7596 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$12590 \$16 \$7029 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12592 \$153 \$7665 \$7632 \$7029 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12593 \$16 \$7029 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12596 \$153 \$7666 \$7632 \$7082 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12597 \$153 \$7634 \$7327 \$7597 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12598 \$153 \$7505 \$7215 \$7388 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12599 \$153 \$7372 \$7550 \$7029 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12600 \$16 \$7709 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12601 \$16 \$7667 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12602 \$16 \$7082 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12604 \$153 \$7389 \$7550 \$7082 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12605 \$16 \$7668 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12606 \$16 \$7130 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12607 \$16 \$7082 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12608 \$153 \$7669 \$7635 \$7082 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12609 \$16 \$8794 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12610 \$153 \$7670 \$7482 \$7571 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12611 \$16 \$7445 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12612 \$16 \$7129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12613 \$16 \$7495 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12616 \$16 \$7387 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12617 \$16 \$6656 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12618 \$16 \$7029 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12619 \$153 \$7671 \$7636 \$7029 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12620 \$153 \$7637 \$6582 \$7613 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12621 \$153 \$7507 \$7327 \$7317 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12622 \$16 \$7540 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12623 \$16 \$7387 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12624 \$153 \$7539 \$7490 \$7317 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12625 \$16 \$7540 \$16 \$153 \$7317 VNB sky130_fd_sc_hd__inv_1
X$12627 \$153 \$7170 \$7686 \$7672 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$12628 \$16 \$7082 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12629 \$153 \$7674 \$7065 \$7726 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12630 \$153 \$7491 \$7171 \$7387 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12631 \$153 \$7598 \$7366 \$7264 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12633 \$16 \$7429 \$7673 \$7599 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$12635 \$16 \$7614 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12636 \$16 \$7129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12637 \$16 \$7129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12638 \$153 \$7687 \$7638 \$7129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12639 \$16 \$7695 \$7673 \$7600 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$12640 \$153 \$7601 \$7638 \$7387 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12641 \$153 \$7601 \$7490 \$7728 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12643 \$16 \$7431 \$16 \$153 \$7417 VNB sky130_fd_sc_hd__inv_1
X$12645 \$153 \$7675 \$7327 \$7728 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12646 \$16 \$7431 \$7673 \$7676 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$12647 \$16 \$7049 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12648 \$153 \$7541 \$7347 \$7574 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$12649 \$153 \$7575 \$7541 \$7307 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12651 \$153 \$7640 \$7639 \$7451 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12653 \$16 \$7641 \$16 \$153 \$7695 VNB sky130_fd_sc_hd__clkbuf_2
X$12654 \$153 \$7640 \$7541 \$7464 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12655 \$153 \$7603 \$7541 \$7131 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12657 \$16 \$7174 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12658 \$153 \$7677 \$7642 \$7174 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12662 \$153 \$7604 \$7375 \$7148 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12664 \$16 \$7133 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12665 \$153 \$7605 \$7643 \$7133 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12666 \$153 \$7678 \$7643 \$7377 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12667 \$153 \$7605 \$7180 \$7734 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12668 \$16 \$8220 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12670 \$16 \$7615 \$16 \$153 \$7049 VNB sky130_fd_sc_hd__clkbuf_2
X$12671 \$153 \$7243 \$8794 \$7509 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$12672 \$153 \$7606 \$7242 \$7464 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12673 \$153 \$7606 \$7639 \$7149 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12674 \$16 \$7668 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12675 \$16 \$7667 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12676 \$153 \$7578 \$7607 \$7392 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12679 \$153 \$7679 \$7180 \$7616 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12680 \$153 \$7644 \$7607 \$7616 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12681 \$16 \$7680 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12683 \$153 \$7645 \$7376 \$7616 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12684 \$153 \$7812 \$7208 \$7616 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12685 \$16 \$7489 \$7496 \$7579 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$12686 \$153 \$7646 \$7639 \$7580 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12689 \$153 \$7681 \$7688 \$7147 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12690 \$153 \$7531 \$7607 \$7580 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12691 \$16 \$7693 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12692 \$16 \$7464 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12693 \$153 \$7617 \$7180 \$7217 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12694 \$153 \$7513 \$7375 \$7318 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12695 \$153 \$7581 \$7639 \$7318 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12697 \$153 \$7428 \$7607 \$7318 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12698 \$153 \$7647 \$7306 \$7582 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$12699 \$153 \$7689 \$7647 \$7464 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12700 \$153 \$5145 \$3719 \$5158 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12701 \$16 \$5158 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12702 \$16 \$5158 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12703 \$16 \$5145 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12704 \$16 \$7147 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12707 \$153 \$7682 \$7497 \$7353 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12708 \$153 \$7312 \$7180 \$7518 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12710 \$153 \$7313 \$7607 \$7518 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12711 \$153 \$7683 \$7497 \$7307 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12712 \$16 \$7307 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12715 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$12716 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$12717 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$12719 \$153 \$7736 \$7544 \$6981 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12720 \$153 \$7648 \$6749 \$7552 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12722 \$16 \$6981 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12723 \$153 \$7618 \$7544 \$6907 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12724 \$16 \$6907 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12726 \$153 \$7553 \$7544 \$6979 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12727 \$153 \$7650 \$6719 \$7552 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12728 \$153 \$7278 \$6913 \$6855 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12730 \$16 \$7545 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12731 \$16 \$7545 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12732 \$153 \$7712 \$6719 \$7711 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12733 \$153 \$7737 \$7784 \$6907 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12734 \$16 \$6907 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12735 \$153 \$7738 \$7620 \$6784 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12736 \$153 \$7738 \$6794 \$7587 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12738 \$16 \$6784 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12739 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$12740 \$153 \$7739 \$7620 \$6783 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12741 \$16 \$6783 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12742 \$16 \$7521 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12743 \$153 \$7740 \$7546 \$6981 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12744 \$153 \$7554 \$6930 \$7140 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12745 \$16 \$6981 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12746 \$16 \$6811 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12747 \$16 \$6733 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12749 \$153 \$7690 \$7546 \$6907 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12750 \$153 \$6811 \$6719 \$6733 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12751 \$16 \$7663 \$16 \$153 \$7608 VNB sky130_fd_sc_hd__inv_1
X$12752 \$16 \$6907 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12753 \$16 \$7466 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12755 \$153 \$7702 \$7701 \$6792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12756 \$16 \$6792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12758 \$16 \$6979 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12759 \$16 \$6883 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12761 \$153 \$7740 \$6930 \$7608 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12762 \$16 \$6784 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12763 \$16 \$6860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12765 \$153 \$7742 \$7703 \$6907 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12766 \$153 \$7556 \$7236 \$6981 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12767 \$153 \$7704 \$6913 \$7609 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12770 \$153 \$7654 \$6749 \$7437 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12771 \$16 \$7713 \$16 \$153 \$6987 VNB sky130_fd_sc_hd__clkbuf_2
X$12772 \$16 \$7714 \$16 \$153 \$6989 VNB sky130_fd_sc_hd__clkbuf_2
X$12773 \$153 \$7622 \$7337 \$6907 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12774 \$16 \$6979 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12776 \$153 \$7771 \$7705 \$7379 \$7785 \$7770 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$12777 \$153 \$7219 \$6913 \$7437 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12778 \$16 \$6907 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12781 \$16 \$7288 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12782 \$153 \$7456 \$7472 \$7623 \$7470 \$7440 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$12783 \$153 \$7472 \$7470 \$7715 \$7456 \$7440 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$12784 \$16 \$7706 \$16 \$153 \$7440 VNB sky130_fd_sc_hd__clkbuf_2
X$12785 \$16 \$7715 \$16 \$153 \$6910 VNB sky130_fd_sc_hd__clkbuf_2
X$12787 \$153 \$7716 \$7006 \$6695 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12788 \$153 \$7743 \$7624 \$6797 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12791 \$16 \$6797 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12792 \$16 \$6991 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12793 \$16 \$7922 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12794 \$153 \$7625 \$7624 \$6754 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12795 \$16 \$6754 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12796 \$16 \$7044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12797 \$153 \$7744 \$7624 \$6771 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12798 \$153 \$7744 \$6865 \$7611 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12799 \$16 \$6771 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12800 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$12802 \$153 \$7628 \$7627 \$7060 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12803 \$16 \$7060 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12804 \$153 \$7629 \$7627 \$6754 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12805 \$153 \$7745 \$7627 \$6797 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12806 \$16 \$6797 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12807 \$16 \$6771 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12810 \$153 \$7717 \$6867 \$7718 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12811 \$153 \$7563 \$6992 \$7043 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12812 \$153 \$7746 \$7707 \$6797 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12813 \$16 \$7466 \$7163 \$7630 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$12815 \$153 \$7747 \$7684 \$6862 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12817 \$153 \$7564 \$6867 \$7043 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12818 \$153 \$7661 \$6324 \$7043 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12820 \$153 \$7534 \$7476 \$7060 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12821 \$153 \$7685 \$6865 \$7458 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12822 \$153 \$7719 \$7006 \$7720 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12823 \$16 \$6771 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12826 \$16 \$7044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12828 \$16 \$6754 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12830 \$16 \$7663 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12831 \$153 \$7721 \$7479 \$6754 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12832 \$153 \$7721 \$6756 \$7612 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12833 \$153 \$7748 \$7479 \$7060 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12834 \$16 \$6991 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12835 \$16 \$7060 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12836 \$16 \$7044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12839 \$153 \$7748 \$6324 \$7612 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12840 \$16 \$7535 \$16 \$153 \$7749 VNB sky130_fd_sc_hd__inv_1
X$12841 \$153 \$7750 \$7708 \$6797 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12842 \$153 \$7750 \$6906 \$7749 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12843 \$16 \$6797 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12845 \$153 \$7751 \$7708 \$6862 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12847 \$153 \$7722 \$6865 \$7749 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12848 \$16 \$6862 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12849 \$16 \$7082 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12850 \$153 \$7752 \$7549 \$7239 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12851 \$16 \$7239 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12852 \$16 \$7067 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12853 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$12854 \$153 \$7631 \$7549 \$7328 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12855 \$16 \$7328 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12858 \$16 \$7387 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12859 \$153 \$7665 \$7066 \$7597 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12860 \$153 \$7753 \$7632 \$7387 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12861 \$153 \$7753 \$7490 \$7597 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12863 \$153 \$7634 \$7632 \$7445 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12864 \$16 \$7709 \$16 \$153 \$7597 VNB sky130_fd_sc_hd__inv_1
X$12866 \$16 \$7328 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12868 \$16 \$7029 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12869 \$16 \$7350 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12871 \$153 \$7723 \$7490 \$7388 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12872 \$153 \$7724 \$7366 \$7388 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12873 \$16 \$7067 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12875 \$16 \$7667 \$16 \$153 \$7388 VNB sky130_fd_sc_hd__inv_1
X$12876 \$153 \$7550 \$7668 \$7754 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$12878 \$153 \$7669 \$7065 \$7571 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12880 \$153 \$7755 \$7635 \$7387 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12881 \$153 \$7537 \$7635 \$7129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12882 \$16 \$7387 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12883 \$153 \$7756 \$7636 \$7387 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12884 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$12885 \$16 \$6656 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12888 \$16 \$7691 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12889 \$16 \$7082 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12890 \$153 \$7692 \$7636 \$7082 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12891 \$153 \$7671 \$7066 \$7613 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12892 \$16 \$7489 \$7673 \$7672 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$12893 \$153 \$7674 \$7790 \$7082 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12894 \$16 \$7387 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12896 \$16 \$7693 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12898 \$153 \$7725 \$7066 \$7726 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12899 \$16 \$7686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12900 \$16 \$7489 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12902 \$153 \$7727 \$7490 \$7726 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12904 \$16 \$7429 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12905 \$16 \$7082 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12906 \$153 \$7694 \$7638 \$7082 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12907 \$16 \$7695 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12908 \$153 \$7694 \$7065 \$7728 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12910 \$153 \$7573 \$7215 \$7417 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12911 \$16 \$7239 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12912 \$16 \$7445 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12913 \$153 \$7675 \$7638 \$7445 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12914 \$16 \$7695 \$16 \$153 \$7728 VNB sky130_fd_sc_hd__inv_1
X$12915 \$16 \$7729 \$16 \$153 \$7429 VNB sky130_fd_sc_hd__clkbuf_2
X$12916 \$153 \$7265 \$7306 \$7676 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$12917 \$16 \$7852 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12918 \$16 \$7730 \$16 \$153 \$7540 VNB sky130_fd_sc_hd__clkbuf_2
X$12920 \$153 \$7757 \$7541 \$7133 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12921 \$16 \$7133 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12923 \$153 \$7696 \$7208 \$7731 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12924 \$153 \$7492 \$7541 \$7353 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12925 \$16 \$7147 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12927 \$153 \$7732 \$7607 \$7731 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12930 \$153 \$7697 \$7639 \$7731 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12931 \$153 \$7697 \$7642 \$7464 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12932 \$153 \$7696 \$7642 \$7131 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12934 \$16 \$7147 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12935 \$16 \$8187 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12936 \$153 \$7678 \$7462 \$7734 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12938 \$153 \$7422 \$7462 \$7097 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12939 \$153 \$7733 \$7463 \$7734 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12940 \$16 \$7353 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12941 \$16 \$7131 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12942 \$153 \$7577 \$7376 \$7734 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12943 \$153 \$7510 \$7462 \$7149 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12944 \$153 \$7758 \$7242 \$7307 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12946 \$16 \$7307 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12948 \$153 \$7735 \$7463 \$7149 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12950 \$16 \$7133 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12951 \$153 \$7679 \$7710 \$7133 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12952 \$16 \$7904 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12953 \$16 \$7667 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12954 \$16 \$7174 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12955 \$153 \$7645 \$7710 \$7174 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12956 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$12959 \$16 \$7464 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12960 \$153 \$7646 \$7688 \$7464 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12961 \$16 \$7489 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12963 \$16 \$7133 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12964 \$16 \$7147 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12965 \$153 \$7759 \$7688 \$7133 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12966 \$153 \$7681 \$7463 \$7580 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12967 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$12968 \$16 \$7147 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12970 \$153 \$7760 \$7698 \$7147 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12972 \$153 \$7699 \$7698 \$7174 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12973 \$153 \$7700 \$7698 \$7464 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12974 \$16 \$7464 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12975 \$16 \$7464 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12977 \$16 \$7174 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12979 \$153 \$7761 \$7647 \$7174 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12980 \$153 \$5534 \$3860 \$5158 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12981 \$16 \$7431 \$16 \$153 \$7782 VNB sky130_fd_sc_hd__inv_1
X$12983 \$153 \$7762 \$7647 \$7147 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12984 \$153 \$7432 \$7375 \$7518 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12985 \$16 \$7464 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12987 \$16 \$7695 \$16 \$153 \$7763 VNB sky130_fd_sc_hd__inv_1
X$12989 \$153 \$7764 \$7497 \$7464 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12990 \$153 \$7211 \$7376 \$7518 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$12991 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$12993 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$12995 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$12996 \$153 \$10997 \$10962 \$10427 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$12997 \$16 \$10427 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$12998 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$13000 \$153 \$10938 \$10962 \$10200 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13001 \$153 \$10938 \$10088 \$11055 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13002 \$16 \$10200 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13005 \$153 \$10904 \$10962 \$10226 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13006 \$153 \$10729 \$10888 \$10842 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$13007 \$16 \$10226 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13009 \$16 \$11078 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13010 \$153 \$10905 \$10963 \$10295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13011 \$16 \$10295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13012 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$13014 \$153 \$10964 \$10161 \$10884 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13015 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$13017 \$153 \$10965 \$10330 \$10884 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13019 \$16 \$10744 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13021 \$16 \$10939 \$10468 \$10998 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$13022 \$16 \$10953 \$16 \$153 \$10468 VNB sky130_fd_sc_hd__clkbuf_2
X$13023 \$16 \$10939 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13025 \$16 \$10890 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13026 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$13028 \$16 \$10295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13030 \$153 \$10999 \$10966 \$10295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13032 \$153 \$10967 \$10161 \$11056 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13033 \$153 \$10940 \$10966 \$10367 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13034 \$153 \$10940 \$10330 \$11056 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13035 \$16 \$10367 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13037 \$16 \$10825 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13040 \$16 \$10367 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13041 \$16 \$9200 \$16 \$153 \$10953 VNB sky130_fd_sc_hd__clkbuf_2
X$13043 \$153 \$10968 \$11000 \$10646 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13044 \$153 \$10968 \$10318 \$10954 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13045 \$153 \$10969 \$10276 \$10954 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13046 \$153 \$10970 \$10705 \$10954 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13047 \$16 \$10476 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13048 \$16 \$10646 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13051 \$153 \$11001 \$10971 \$10368 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13052 \$153 \$11029 \$10330 \$11057 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13053 \$16 \$10368 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13054 \$153 \$11002 \$10817 \$10476 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13055 \$153 \$11002 \$10705 \$10805 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13056 \$16 \$10646 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13057 \$16 \$10226 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13059 \$153 \$11003 \$10817 \$10200 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13060 \$153 \$11181 \$10817 \$10295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13061 \$153 \$10886 \$10885 \$10878 \$10877 \$10907 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$13062 \$153 \$10885 \$10907 \$10955 \$10877 \$10878 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$13063 \$16 \$10955 \$16 \$153 \$10764 VNB sky130_fd_sc_hd__clkbuf_2
X$13066 \$16 \$10764 \$10525 \$10908 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$13067 \$16 \$11004 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13068 \$16 \$11078 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13069 \$153 \$10909 \$10821 \$10514 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13070 \$16 \$11078 \$16 \$153 \$10941 VNB sky130_fd_sc_hd__inv_1
X$13071 \$153 \$10910 \$10516 \$10941 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13072 \$153 \$10769 \$10344 \$10941 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13073 \$153 \$10770 \$10686 \$10477 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13076 \$153 \$10889 \$10821 \$10382 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13078 \$153 \$10942 \$10822 \$10526 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13079 \$153 \$11005 \$10822 \$10514 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13080 \$16 \$10526 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13081 \$16 \$10744 \$10525 \$10943 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$13083 \$153 \$10942 \$10516 \$10750 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13084 \$153 \$11033 \$10686 \$10750 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13085 \$153 \$10972 \$10247 \$10956 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13086 \$153 \$11034 \$10516 \$10956 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13087 \$153 \$10773 \$10344 \$10647 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13088 \$16 \$11993 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13089 \$153 \$10911 \$10686 \$10647 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13091 \$153 \$10973 \$10098 \$10956 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13092 \$16 \$9550 \$16 \$153 \$11123 VNB sky130_fd_sc_hd__clkbuf_2
X$13093 \$16 \$9550 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13094 \$153 \$10752 \$10731 \$10606 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13095 \$153 \$10912 \$10309 \$10891 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13096 \$16 \$10606 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13097 \$16 \$10825 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13099 \$153 \$10957 \$10401 \$10958 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13102 \$16 \$10470 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13103 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$13105 \$153 \$11006 \$11049 \$10606 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13106 \$16 \$10606 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13107 \$16 \$10413 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13109 \$16 \$10605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13111 \$153 \$10914 \$10893 \$10470 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13113 \$153 \$10915 \$10516 \$10892 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13114 \$16 \$10974 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13115 \$16 \$10959 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13116 \$153 \$10944 \$10893 \$10298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13117 \$153 \$10944 \$10401 \$10892 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13118 \$16 \$10298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13119 \$153 \$10945 \$10975 \$10382 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13121 \$153 \$11007 \$10975 \$10514 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13122 \$153 \$10896 \$10975 \$10338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13123 \$153 \$11008 \$10975 \$10470 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13124 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$13125 \$16 \$10473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13127 \$153 \$10895 \$10733 \$10473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13128 \$153 \$10808 \$10733 \$10551 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13129 \$16 \$10551 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13131 \$16 \$10831 \$11127 \$10917 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$13132 \$153 \$10980 \$10734 \$10386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13134 \$153 \$10976 \$10472 \$11207 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13135 \$153 \$10846 \$10833 \$10609 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13136 \$16 \$11207 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13137 \$16 \$10831 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13139 \$153 \$10977 \$10471 \$10480 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13140 \$16 \$10978 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13141 \$16 \$10386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13142 \$153 \$11009 \$10979 \$10386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13143 \$16 \$10854 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13144 \$16 \$10739 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13146 \$153 \$10980 \$10472 \$10480 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13147 \$153 \$11091 \$10919 \$10810 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13148 \$153 \$11146 \$10714 \$10810 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13149 \$153 \$11010 \$10881 \$10551 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13151 \$153 \$11041 \$10501 \$10946 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13152 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$13154 \$153 \$10920 \$10919 \$10946 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13155 \$153 \$11011 \$10882 \$10386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13156 \$153 \$10871 \$10417 \$10811 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13158 \$16 \$10473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13159 \$16 \$10386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13160 \$153 \$10882 \$10981 \$10921 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$13161 \$16 \$10661 \$16 \$153 \$10811 VNB sky130_fd_sc_hd__inv_1
X$13163 \$153 \$11011 \$10472 \$10811 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13164 \$16 \$10552 \$16 \$153 \$10757 VNB sky130_fd_sc_hd__inv_1
X$13166 \$153 \$10947 \$10834 \$10386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13167 \$153 \$10982 \$10417 \$10923 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13168 \$153 \$10947 \$10472 \$10923 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13169 \$153 \$10983 \$10833 \$10948 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13171 \$16 \$10649 \$16 \$153 \$10923 VNB sky130_fd_sc_hd__inv_1
X$13172 \$16 \$10473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13173 \$16 \$10473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13174 \$153 \$10984 \$10919 \$10923 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13175 \$153 \$10924 \$10501 \$10923 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13176 \$16 \$10386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13177 \$153 \$10949 \$10658 \$10473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13178 \$153 \$10949 \$10501 \$10926 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13179 \$16 \$10853 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13180 \$16 \$10409 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13182 \$16 \$10960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13183 \$153 \$10658 \$10960 \$10985 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$13184 \$16 \$10409 \$10737 \$10985 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$13185 \$16 \$10860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13187 \$153 \$10927 \$10417 \$10926 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13189 \$16 \$10986 \$16 \$153 \$10987 VNB sky130_fd_sc_hd__clkbuf_2
X$13190 \$16 \$11253 \$16 \$153 \$11012 VNB sky130_fd_sc_hd__clkbuf_2
X$13191 \$153 \$10898 \$10950 \$10988 \$11012 \$10987 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$13192 \$16 \$11147 \$16 \$153 \$10950 VNB sky130_fd_sc_hd__clkbuf_2
X$13194 \$153 \$10899 \$10950 \$11012 \$10987 \$10988 \$16 \$16 VNB
+ sky130_fd_sc_hd__nor4b_2
X$13195 \$153 \$10950 \$10987 \$10900 \$11012 \$10988 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$13196 \$16 \$10989 \$16 \$153 \$11013 VNB sky130_fd_sc_hd__clkbuf_2
X$13197 \$153 \$11014 \$10839 \$10392 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13198 \$153 \$10930 \$10642 \$10812 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13199 \$16 \$10392 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13200 \$16 \$11015 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13201 \$16 \$11016 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13203 \$16 \$10831 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13204 \$153 \$10931 \$10587 \$10812 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13205 \$153 \$10951 \$10839 \$10617 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13206 \$153 \$10951 \$10560 \$10812 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13207 \$16 \$10617 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13209 \$153 \$11017 \$11052 \$10617 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13212 \$153 \$11017 \$10560 \$10961 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13213 \$153 \$10790 \$10815 \$10518 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13214 \$16 \$10990 \$16 \$153 \$10838 VNB sky130_fd_sc_hd__clkbuf_2
X$13215 \$16 \$9550 \$16 \$153 \$10990 VNB sky130_fd_sc_hd__clkbuf_2
X$13216 \$153 \$10991 \$10560 \$10814 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13217 \$153 \$10992 \$10285 \$10814 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13218 \$153 \$10993 \$10587 \$10814 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13220 \$16 \$10552 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13223 \$153 \$10952 \$10901 \$10346 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13224 \$153 \$10952 \$10285 \$10902 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13225 \$16 \$10552 \$10644 \$11018 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$13226 \$153 \$10994 \$10560 \$10902 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13227 \$153 \$11019 \$10995 \$10467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13230 \$153 \$10859 \$10560 \$10858 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13231 \$153 \$11020 \$10995 \$10446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13232 \$16 \$10981 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13234 \$16 \$10661 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13235 \$16 \$10393 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13236 \$153 \$11021 \$10995 \$10393 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13237 \$16 \$10852 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13238 \$16 \$10853 \$10644 \$10996 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$13240 \$16 \$10597 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13241 \$16 \$10860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13242 \$153 \$10796 \$10852 \$10996 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$13243 \$16 \$10853 \$16 \$153 \$11022 VNB sky130_fd_sc_hd__inv_1
X$13244 \$153 \$10422 \$10694 \$10521 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13245 \$153 \$9782 \$9122 \$10222 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13246 \$153 \$9919 \$9103 \$10222 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13247 \$16 \$10222 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13248 \$16 \$10393 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13249 \$16 \$10393 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13250 \$16 \$10346 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13252 \$16 \$10529 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13253 \$16 \$10853 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13254 \$16 \$10326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13255 \$153 \$11023 \$10796 \$10326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13256 \$16 \$10510 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13258 \$16 \$10510 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13259 \$153 \$11024 \$10796 \$10446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13261 \$16 \$7033 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13262 \$153 \$8086 \$7462 \$7033 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13264 \$16 \$8086 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13265 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$13266 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$13267 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$13269 \$153 \$11070 \$10962 \$10368 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13270 \$16 \$10368 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13271 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$13273 \$153 \$11070 \$10303 \$11055 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13274 \$153 \$11048 \$10276 \$11055 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13276 \$153 \$10903 \$10330 \$10511 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13277 \$153 \$11025 \$10962 \$10476 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13278 \$153 \$11025 \$10705 \$11055 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13279 \$16 \$11078 \$16 \$153 \$11055 VNB sky130_fd_sc_hd__inv_1
X$13281 \$16 \$11078 \$10468 \$11072 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$13283 \$153 \$11026 \$10963 \$10646 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13284 \$153 \$11026 \$10318 \$10884 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13285 \$16 \$10646 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13287 \$153 \$11073 \$10963 \$10368 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13288 \$16 \$10368 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13289 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$13291 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$13292 \$153 \$11074 \$10532 \$10200 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13293 \$16 \$10939 \$16 \$153 \$10745 VNB sky130_fd_sc_hd__inv_1
X$13294 \$16 \$10200 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13295 \$16 \$10939 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13296 \$153 \$11027 \$10966 \$10646 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13298 \$153 \$11027 \$10318 \$11056 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13299 \$16 \$10226 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13302 \$153 \$10999 \$10276 \$11056 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13304 \$16 \$10427 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13305 \$153 \$11028 \$10966 \$10427 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13306 \$153 \$11076 \$10966 \$10476 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13307 \$153 \$11028 \$10327 \$11056 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13308 \$16 \$10476 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13311 \$153 \$10970 \$11000 \$10476 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13312 \$16 \$10476 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13313 \$16 \$11993 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13315 \$16 \$10367 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13316 \$153 \$11029 \$10971 \$10367 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13317 \$153 \$11001 \$10303 \$11057 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13318 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$13319 \$16 \$10624 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13320 \$16 \$10427 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13322 \$153 \$11030 \$10817 \$10427 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13323 \$153 \$11030 \$10327 \$10805 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13324 \$153 \$11031 \$10817 \$10368 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13325 \$153 \$11031 \$10303 \$10805 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13326 \$16 \$10368 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13327 \$16 \$11058 \$16 \$153 \$11078 VNB sky130_fd_sc_hd__clkbuf_2
X$13330 \$153 \$10820 \$10877 \$10878 \$10885 \$10907 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$13331 \$153 \$10877 \$10885 \$11079 \$10907 \$10878 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$13332 \$16 \$10865 \$16 \$153 \$10744 VNB sky130_fd_sc_hd__clkbuf_2
X$13333 \$16 \$6667 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13334 \$153 \$10821 \$11004 \$11080 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$13335 \$153 \$11081 \$10821 \$10605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13337 \$16 \$10514 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13338 \$153 \$11082 \$10821 \$10338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13339 \$16 \$10764 \$16 \$153 \$10750 VNB sky130_fd_sc_hd__inv_1
X$13341 \$153 \$11032 \$10821 \$10298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13342 \$153 \$11032 \$10401 \$10941 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13343 \$153 \$11059 \$10247 \$10941 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13345 \$16 \$10382 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13346 \$153 \$11033 \$10822 \$10605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13347 \$16 \$10605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13348 \$16 \$10514 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13349 \$16 \$10939 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13350 \$16 \$11114 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13351 \$153 \$11060 \$11114 \$11083 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$13352 \$153 \$11034 \$11060 \$10526 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13354 \$16 \$10526 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13355 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$13356 \$153 \$11035 \$11060 \$10298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13357 \$153 \$11035 \$10401 \$10956 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13358 \$16 \$10298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13360 \$153 \$11036 \$11124 \$10606 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13361 \$16 \$10606 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13362 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$13364 \$153 \$11037 \$11124 \$10338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13365 \$153 \$11037 \$10309 \$10958 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13367 \$153 \$11038 \$11049 \$10514 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13368 \$153 \$11038 \$10538 \$11061 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13369 \$16 \$10514 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13371 \$16 \$10706 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13373 \$153 \$10893 \$10706 \$10913 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$13374 \$153 \$11006 \$10344 \$11061 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13376 \$16 \$10413 \$16 \$153 \$10892 VNB sky130_fd_sc_hd__inv_1
X$13377 \$16 \$10470 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13378 \$16 \$10413 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13379 \$153 \$11062 \$10309 \$10892 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13380 \$153 \$11085 \$10893 \$10605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13382 \$153 \$10916 \$10098 \$10892 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13384 \$16 \$10298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13385 \$153 \$11087 \$10975 \$10298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13386 \$16 \$10514 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13387 \$16 \$10974 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13389 \$153 \$11007 \$10538 \$10894 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13390 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$13391 \$16 \$10526 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13392 \$153 \$11008 \$10247 \$10894 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13395 \$16 \$10470 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13397 \$153 \$11063 \$10516 \$10894 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13398 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$13399 \$16 \$10809 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13400 \$153 \$11088 \$11050 \$10809 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13401 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$13402 \$153 \$11089 \$11050 \$10611 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13404 \$153 \$11064 \$10501 \$11209 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13405 \$153 \$11089 \$10833 \$11209 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13406 \$153 \$11039 \$10734 \$10735 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13407 \$153 \$11039 \$10919 \$10480 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13408 \$153 \$11090 \$10472 \$11065 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13409 \$16 \$10978 \$16 \$153 \$10480 VNB sky130_fd_sc_hd__inv_1
X$13413 \$16 \$10809 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13414 \$16 \$11015 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13416 \$16 \$10735 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13417 \$153 \$11091 \$10979 \$10735 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13418 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$13420 \$16 \$10578 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13421 \$153 \$11040 \$10979 \$10578 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13422 \$153 \$11040 \$10370 \$10810 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13424 \$153 \$11041 \$10881 \$10473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13425 \$153 \$11010 \$10471 \$10946 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13426 \$153 \$10848 \$10833 \$10946 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13428 \$16 \$10386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13429 \$153 \$11042 \$10882 \$10611 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13431 \$16 \$10981 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13433 \$153 \$11094 \$10471 \$10811 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13434 \$16 \$11212 \$16 \$153 \$10737 VNB sky130_fd_sc_hd__clkbuf_2
X$13435 \$16 \$10735 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13436 \$153 \$11043 \$10882 \$10735 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13437 \$153 \$11043 \$10919 \$10811 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13438 \$153 \$10982 \$10834 \$10300 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13441 \$16 \$10649 \$10737 \$11051 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$13442 \$153 \$10834 \$12050 \$11051 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$13443 \$153 \$11044 \$10834 \$10551 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13444 \$153 \$11044 \$10471 \$10923 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13445 \$153 \$10785 \$10833 \$10517 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13446 \$16 \$10578 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13448 \$153 \$11096 \$11066 \$10578 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13449 \$16 \$10735 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13450 \$153 \$11067 \$11066 \$10735 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13451 \$16 \$10300 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13452 \$16 \$10809 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13453 \$153 \$11098 \$11066 \$10809 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13454 \$16 \$6540 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13456 \$153 \$11067 \$10919 \$11099 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13457 \$16 \$6540 \$16 \$153 \$10986 VNB sky130_fd_sc_hd__clkbuf_2
X$13458 \$153 \$10835 \$11012 \$10988 \$10950 \$10987 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$13459 \$153 \$10836 \$10987 \$10988 \$11012 \$10950 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$13460 \$153 \$11012 \$10950 \$10928 \$10987 \$10988 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$13461 \$16 \$10978 \$10838 \$11100 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$13462 \$153 \$11068 \$10815 \$11016 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13464 \$153 \$10839 \$11015 \$11100 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$13465 \$16 \$11069 \$16 \$153 \$10552 VNB sky130_fd_sc_hd__clkbuf_2
X$13466 \$16 \$10392 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13467 \$153 \$11045 \$11052 \$10326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13468 \$153 \$11045 \$10466 \$10961 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13469 \$16 \$10326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13470 \$153 \$10932 \$10376 \$10812 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13472 \$153 \$11101 \$10587 \$10961 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13473 \$153 \$11046 \$11052 \$10346 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13474 \$153 \$11046 \$10285 \$10961 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13475 \$16 \$10346 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13476 \$153 \$10992 \$10740 \$10346 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13477 \$16 \$10346 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13478 \$16 \$11013 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13480 \$16 \$10564 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13481 \$153 \$11104 \$10740 \$10564 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13482 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$13483 \$16 \$10393 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13484 \$153 \$11047 \$10901 \$10393 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13485 \$153 \$11047 \$10694 \$10902 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13486 \$16 \$10346 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13487 \$16 \$10617 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13488 \$16 \$10990 \$16 \$153 \$10644 VNB sky130_fd_sc_hd__clkbuf_2
X$13490 \$153 \$10994 \$10901 \$10617 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13491 \$16 \$10467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13492 \$16 \$10564 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13493 \$153 \$11105 \$10995 \$10564 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13494 \$153 \$11106 \$10995 \$10346 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13495 \$16 \$10346 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13498 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$13499 \$16 \$10617 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13500 \$153 \$11107 \$10995 \$10617 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13501 \$153 \$10566 \$10694 \$10650 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13502 \$153 \$10421 \$10285 \$10650 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13504 \$153 \$11108 \$11053 \$10393 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13506 \$153 \$10450 \$10466 \$10521 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13507 \$153 \$11109 \$11053 \$10346 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13508 \$153 \$10631 \$10642 \$10521 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13509 \$153 \$10423 \$10285 \$10521 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13511 \$153 \$10632 \$10642 \$10741 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13512 \$16 \$10446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13514 \$16 \$10617 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13515 \$153 \$11110 \$10796 \$10467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13516 \$16 \$10510 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13517 \$16 \$10510 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13518 \$153 \$11054 \$8977 \$10510 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13519 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$13520 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$13521 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$13522 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$13523 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$13524 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$13525 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$13526 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$13528 \$153 \$12716 \$12412 \$12512 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13529 \$153 \$12638 \$12656 \$12294 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13531 \$153 \$12790 \$12656 \$12152 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13532 \$153 \$12716 \$12656 \$12230 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13534 \$153 \$12685 \$12656 \$12158 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13535 \$16 \$12294 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13536 \$16 \$12152 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13538 \$16 \$12230 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13539 \$153 \$12685 \$12057 \$12512 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13540 \$153 \$12655 \$12134 \$12512 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13541 \$16 \$12158 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13542 \$153 \$12585 \$12656 \$12095 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13543 \$16 \$11636 \$12779 \$12791 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$13544 \$153 \$12717 \$12229 \$12512 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13546 \$153 \$12513 \$12656 \$12003 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13547 \$153 \$12717 \$12656 \$12093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13548 \$16 \$12003 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13550 \$153 \$12754 \$12469 \$12294 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13551 \$153 \$12754 \$12208 \$12563 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13553 \$16 \$12093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13555 \$16 \$11369 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13556 \$16 \$12236 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13557 \$16 \$12294 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13558 \$16 \$11369 \$12779 \$12792 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$13560 \$153 \$12614 \$12469 \$12152 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13561 \$153 \$12793 \$12469 \$12230 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13563 \$153 \$12707 \$12209 \$12426 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13566 \$16 \$12564 \$16 \$153 \$12779 VNB sky130_fd_sc_hd__clkbuf_2
X$13567 \$153 \$12707 \$12586 \$12152 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13568 \$153 \$12639 \$12586 \$12294 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13569 \$16 \$12152 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13570 \$16 \$12294 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13571 \$16 \$12236 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13572 \$16 \$11190 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13573 \$16 \$10939 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13574 \$16 \$11567 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13578 \$153 \$12718 \$12586 \$12158 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13579 \$153 \$12640 \$12586 \$12230 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13580 \$16 \$12158 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13581 \$153 \$12718 \$12057 \$12426 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13582 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$13583 \$153 \$12719 \$12471 \$12152 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13584 \$16 \$12230 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13587 \$153 \$12470 \$11810 \$12578 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13588 \$153 \$12719 \$12209 \$12578 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13589 \$153 \$12657 \$12208 \$12578 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13590 \$16 \$12158 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13592 \$16 \$12152 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13593 \$16 \$11297 \$12015 \$12701 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$13594 \$153 \$12794 \$12720 \$12095 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13596 \$153 \$12720 \$11364 \$12701 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$13597 \$16 \$11297 \$16 \$153 \$12780 VNB sky130_fd_sc_hd__inv_1
X$13598 \$16 \$12095 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13599 \$153 \$12658 \$12412 \$12578 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13600 \$16 \$11364 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13602 \$153 \$12721 \$12444 \$12294 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13603 \$16 \$11297 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13606 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$13608 \$153 \$12721 \$12208 \$12413 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13609 \$153 \$12722 \$12444 \$12152 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13610 \$153 \$12763 \$12444 \$12230 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13611 \$16 \$12294 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13612 \$16 \$12152 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13615 \$153 \$12589 \$12057 \$12413 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13616 \$153 \$12763 \$12412 \$12413 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13617 \$16 \$12230 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13618 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$13620 \$153 \$12796 \$12514 \$12230 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13621 \$153 \$12723 \$12514 \$12152 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13623 \$16 \$12230 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13624 \$16 \$12152 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13627 \$153 \$12723 \$12209 \$12579 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13628 \$153 \$12724 \$12514 \$12294 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13629 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$13630 \$153 \$12724 \$12208 \$12579 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13631 \$16 \$11594 \$12897 \$12913 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$13632 \$153 \$12702 \$12391 \$12230 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13633 \$16 \$12294 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13635 \$16 \$11594 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13637 \$153 \$12702 \$12412 \$12392 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13638 \$153 \$12797 \$12708 \$12003 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13639 \$153 \$12725 \$12391 \$12152 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13641 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$13642 \$16 \$12003 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13644 \$153 \$12726 \$12708 \$12093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13645 \$153 \$12727 \$12708 \$12236 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13646 \$16 \$12093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13647 \$153 \$12726 \$12229 \$12783 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13649 \$16 \$11078 \$12159 \$12661 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$13651 \$16 \$12236 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13652 \$153 \$12727 \$12134 \$12783 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13653 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$13655 \$153 \$12728 \$12615 \$12044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13657 \$153 \$12755 \$12615 \$12259 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13658 \$16 \$12044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13661 \$153 \$12755 \$12307 \$12641 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13662 \$153 \$12756 \$12615 \$12295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13663 \$153 \$12728 \$12068 \$12641 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13664 \$153 \$12757 \$12615 \$12083 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13665 \$153 \$12756 \$12155 \$12641 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13668 \$16 \$11078 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13669 \$16 \$12160 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13670 \$16 \$12083 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13671 \$153 \$12709 \$12615 \$12101 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13673 \$153 \$12757 \$12174 \$12641 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13674 \$153 \$12709 \$12476 \$12641 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13675 \$16 \$12101 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13676 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$13677 \$16 \$12101 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13678 \$16 \$12101 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13681 \$153 \$12593 \$12068 \$12154 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13682 \$153 \$12686 \$12533 \$12296 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13684 \$153 \$12784 \$12476 \$12781 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13685 \$153 \$12686 \$12359 \$12154 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13686 \$153 \$12662 \$12476 \$12154 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13687 \$16 \$12296 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13689 \$16 \$10523 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13690 \$16 \$11369 \$16 \$153 \$12781 VNB sky130_fd_sc_hd__inv_1
X$13692 \$153 \$12687 \$12477 \$12259 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13693 \$16 \$12044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13694 \$16 \$11369 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13695 \$153 \$12619 \$12477 \$12044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13696 \$153 \$12687 \$12307 \$12498 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13697 \$16 \$12259 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13698 \$16 \$12044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13701 \$16 \$10453 \$16 \$153 \$12729 VNB sky130_fd_sc_hd__inv_1
X$13702 \$153 \$12764 \$12477 \$12296 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13703 \$16 \$10453 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13705 \$153 \$12730 \$12710 \$12083 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13706 \$16 \$12296 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13708 \$153 \$12730 \$12174 \$12729 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13709 \$16 \$12083 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13710 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$13712 \$153 \$12643 \$12710 \$12101 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13714 \$153 \$12765 \$11364 \$12663 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$13715 \$153 \$12644 \$12500 \$12296 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13716 \$16 \$12101 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13717 \$16 \$11297 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13718 \$16 \$11297 \$16 \$153 \$12758 VNB sky130_fd_sc_hd__inv_1
X$13719 \$16 \$12581 \$16 \$153 \$12785 VNB sky130_fd_sc_hd__clkbuf_2
X$13722 \$153 \$12766 \$12765 \$12160 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13723 \$153 \$12731 \$12500 \$12241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13724 \$16 \$12160 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13726 \$16 \$12296 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13727 \$153 \$12767 \$12765 \$12241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13728 \$16 \$12241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13729 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$13732 \$153 \$12664 \$12307 \$12360 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13733 \$153 \$12767 \$12363 \$12758 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13734 \$16 \$12241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13735 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$13737 \$153 \$12731 \$12363 \$12360 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13738 \$153 \$12732 \$12508 \$12296 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13741 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$13742 \$153 \$12732 \$12359 \$12429 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13743 \$153 \$12733 \$12508 \$12241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13744 \$153 \$12798 \$12502 \$12083 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13745 \$16 \$12241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13747 \$16 \$12083 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13749 \$153 \$12703 \$12476 \$12429 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13750 \$153 \$12768 \$12502 \$12160 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13752 \$153 \$12688 \$12502 \$12044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13753 \$153 \$12798 \$12174 \$12430 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13755 \$153 \$12734 \$12502 \$12241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13756 \$16 \$12044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13758 \$16 \$11594 \$12785 \$12915 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$13760 \$153 \$12759 \$12621 \$12259 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13761 \$153 \$12688 \$12068 \$12430 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13763 \$153 \$12769 \$12621 \$12101 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13764 \$16 \$10974 \$16 \$153 \$12704 VNB sky130_fd_sc_hd__inv_1
X$13767 \$153 \$12759 \$12307 \$12704 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13768 \$16 \$12259 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13769 \$153 \$12769 \$12476 \$12704 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13770 \$16 \$12101 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13771 \$16 \$12241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13772 \$16 \$12296 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13773 \$153 \$12735 \$12621 \$12296 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13774 \$153 \$12666 \$12155 \$12704 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13776 \$16 \$11594 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13778 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$13779 \$153 \$12735 \$12359 \$12704 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13781 \$153 \$12399 \$12711 \$12571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13783 \$16 \$12164 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13784 \$16 \$12571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13785 \$153 \$12799 \$12711 \$12164 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13787 \$153 \$12689 \$12711 \$12297 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13788 \$153 \$12770 \$12363 \$12881 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13789 \$153 \$12799 \$12217 \$12690 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13790 \$153 \$12597 \$12309 \$12325 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13791 \$153 \$12689 \$12582 \$12690 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13793 \$16 \$12233 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13795 \$153 \$12771 \$12711 \$12233 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13796 \$16 \$10831 \$16 \$153 \$12690 VNB sky130_fd_sc_hd__inv_1
X$13797 \$153 \$12711 \$12406 \$12668 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$13798 \$153 \$12771 \$12603 \$12690 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13799 \$16 \$12297 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13801 \$16 \$12233 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13803 \$16 \$12297 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13805 \$153 \$12646 \$12482 \$12233 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13807 \$16 \$12326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13808 \$153 \$12772 \$12736 \$12115 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13809 \$153 \$12691 \$12736 \$12326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13810 \$153 \$12772 \$12234 \$12787 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13812 \$153 \$12786 \$12603 \$12787 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13813 \$153 \$12691 \$12264 \$12787 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13814 \$16 \$12164 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13815 \$16 \$12571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13817 \$153 \$12736 \$10780 \$12712 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$13818 \$153 \$12800 \$12736 \$12571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13820 \$16 \$10854 \$12379 \$12712 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$13821 \$16 \$10854 \$16 \$153 \$12787 VNB sky130_fd_sc_hd__inv_1
X$13823 \$153 \$12483 \$12518 \$12571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13824 \$153 \$12647 \$12518 \$12297 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13825 \$16 \$12297 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13826 \$16 \$12571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13828 \$16 \$10854 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13829 \$16 \$12233 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13831 \$16 \$12298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13832 \$153 \$12692 \$12518 \$12233 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13834 \$153 \$12625 \$12518 \$12298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13835 \$153 \$12692 \$12603 \$12503 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13837 \$16 \$11502 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13838 \$16 \$11604 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13839 \$16 \$12298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13840 \$16 \$11622 \$12634 \$12713 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$13841 \$153 \$12773 \$12452 \$12298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13843 \$153 \$12452 \$12612 \$12713 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$13844 \$153 \$12773 \$12165 \$12432 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13846 \$153 \$12649 \$12452 \$12219 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13847 \$16 \$11216 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13848 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$13849 \$16 \$12297 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13851 \$153 \$12760 \$12452 \$12297 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13852 \$153 \$12737 \$12452 \$12233 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13853 \$153 \$12693 \$12670 \$12115 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13854 \$153 \$12760 \$12582 \$12432 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13856 \$153 \$12484 \$12309 \$12200 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13857 \$16 \$12115 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13858 \$16 \$12298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13859 \$153 \$12705 \$12670 \$12298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13860 \$153 \$12693 \$12234 \$12671 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13862 \$153 \$12738 \$12670 \$12297 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13863 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$13865 \$16 \$11496 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13866 \$16 \$11585 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13867 \$153 \$12738 \$12582 \$12671 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13868 \$153 \$12739 \$12670 \$12233 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13869 \$16 \$12233 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13870 \$16 \$12115 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13871 \$153 \$12740 \$12714 \$12115 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13872 \$16 \$10552 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13873 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$13875 \$153 \$12705 \$12165 \$12671 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13876 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$13877 \$153 \$12714 \$12404 \$12801 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$13878 \$153 \$12740 \$12234 \$12706 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13879 \$153 \$12741 \$12714 \$12326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13880 \$16 \$12297 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13881 \$16 \$12326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13882 \$16 \$12404 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13884 \$16 \$12298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13885 \$16 \$11413 \$16 \$153 \$12706 VNB sky130_fd_sc_hd__inv_1
X$13886 \$153 \$12694 \$12714 \$12571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13887 \$153 \$12674 \$12165 \$12488 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13888 \$153 \$12802 \$12605 \$12219 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13889 \$16 \$12571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13890 \$16 \$12164 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13891 \$16 \$12115 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13893 \$153 \$12672 \$12165 \$12333 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13894 \$153 \$12774 \$12605 \$12297 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13895 \$16 \$12298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13896 \$153 \$12742 \$12605 \$12164 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13898 \$153 \$12742 \$12217 \$12488 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13900 \$153 \$12695 \$12605 \$12115 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13902 \$153 \$12775 \$12605 \$12326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13903 \$153 \$12695 \$12234 \$12488 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13904 \$153 \$12775 \$12264 \$12488 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13905 \$16 \$12433 \$12162 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$13906 \$16 \$12433 \$11216 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$13909 \$16 \$12433 \$11842 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$13910 \$16 \$12299 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13911 \$153 \$12803 \$12675 \$12299 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13912 \$153 \$12696 \$12675 \$11983 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13913 \$153 \$12776 \$11942 \$12650 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13915 \$153 \$12696 \$11881 \$12650 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13917 \$16 \$10854 \$16 \$153 \$12650 VNB sky130_fd_sc_hd__inv_1
X$13918 \$16 \$10780 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13920 \$16 \$12303 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13921 \$153 \$12651 \$12675 \$12351 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13922 \$153 \$12743 \$12675 \$12303 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13923 \$153 \$12743 \$12227 \$12650 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13924 \$16 \$12351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13925 \$16 \$10854 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13926 \$16 \$12406 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13930 \$153 \$12715 \$12406 \$12676 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$13931 \$16 \$12303 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13932 \$153 \$12744 \$12715 \$12303 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13933 \$16 \$12120 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13934 \$153 \$12744 \$12227 \$12824 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13936 \$16 \$12010 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13937 \$153 \$12697 \$12715 \$12010 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13938 \$16 \$12287 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13940 \$153 \$12745 \$12715 \$12287 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13941 \$153 \$12697 \$11942 \$12824 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13942 \$16 \$11604 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13943 \$153 \$12745 \$12339 \$12824 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13944 \$16 \$12303 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13945 \$16 \$12299 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13946 \$153 \$12761 \$12489 \$12303 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13948 \$153 \$12746 \$12489 \$12299 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13950 \$153 \$12746 \$12371 \$12337 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13951 \$153 \$12748 \$12489 \$11983 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13952 \$16 \$11983 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13953 \$16 \$11622 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13954 \$16 \$12574 \$16 \$153 \$12747 VNB sky130_fd_sc_hd__clkbuf_2
X$13956 \$153 \$12748 \$11881 \$12337 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13957 \$16 \$11622 \$12747 \$12677 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$13958 \$16 \$12303 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13960 \$153 \$12653 \$12583 \$12351 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13961 \$153 \$12652 \$12583 \$12303 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13962 \$16 \$12351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13965 \$16 \$12299 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13966 \$16 \$11983 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13967 \$153 \$12777 \$12583 \$11983 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13968 \$153 \$12698 \$12583 \$12299 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13969 \$153 \$12698 \$12371 \$12435 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13970 \$153 \$12777 \$11881 \$12435 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13973 \$16 \$12299 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13975 \$16 \$12287 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13976 \$153 \$12699 \$12635 \$12299 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13977 \$153 \$12804 \$12635 \$12287 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13978 \$153 \$12226 \$12119 \$12147 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13980 \$16 \$12404 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13981 \$16 \$12303 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13982 \$153 \$12805 \$12635 \$12303 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13985 \$153 \$12699 \$12371 \$12680 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13986 \$16 \$12120 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13987 \$153 \$12807 \$12404 \$12806 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$13988 \$153 \$12749 \$12635 \$12120 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13990 \$16 \$12384 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$13991 \$153 \$12749 \$12182 \$12680 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13993 \$153 \$12788 \$11942 \$12680 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13995 \$16 \$11413 \$16 \$153 \$12750 VNB sky130_fd_sc_hd__inv_1
X$13996 \$153 \$12681 \$11881 \$12680 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$13997 \$153 \$12611 \$12409 \$11983 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$13998 \$153 \$12808 \$12807 \$11983 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14001 \$153 \$12682 \$12182 \$12521 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14002 \$16 \$12120 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14004 \$16 \$11546 \$12678 \$12778 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$14005 \$153 \$12751 \$12409 \$12287 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14006 \$153 \$12636 \$11385 \$12778 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$14007 \$16 \$12287 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14009 \$16 \$11798 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14010 \$153 \$12751 \$12339 \$12521 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14011 \$16 \$12120 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14012 \$153 \$12752 \$12636 \$12120 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14013 \$153 \$11321 \$10642 \$11322 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14014 \$153 \$11108 \$10694 \$11322 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14015 \$16 \$11546 \$16 \$153 \$12654 VNB sky130_fd_sc_hd__inv_1
X$14016 \$16 \$12287 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14018 \$16 \$12010 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14019 \$153 \$11109 \$10285 \$11322 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14021 \$153 \$12753 \$12636 \$12010 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14022 \$153 \$11174 \$10815 \$11322 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14024 \$153 \$12753 \$11942 \$12654 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14025 \$16 \$12303 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14026 \$153 \$12700 \$12636 \$12303 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14027 \$16 \$12351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14029 \$16 \$12782 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14031 \$16 \$12303 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14032 \$153 \$12633 \$12179 \$12654 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14033 \$153 \$11986 \$10815 \$11926 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14034 \$153 \$12789 \$12119 \$12654 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14035 \$153 \$12700 \$12227 \$12654 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14036 \$153 \$11613 \$10560 \$12782 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14037 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$14039 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$14041 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$14042 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$14043 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$14044 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$14045 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$14046 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$14048 \$153 \$12151 \$12134 \$12150 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14049 \$153 \$12340 \$12209 \$12150 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14050 \$153 \$12183 \$12019 \$12294 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14051 \$153 \$12184 \$12209 \$12020 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14054 \$153 \$12183 \$12208 \$12020 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14055 \$153 \$12184 \$12019 \$12152 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14056 \$153 \$12090 \$12057 \$12020 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14057 \$153 \$12250 \$12019 \$12236 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14058 \$16 \$12294 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14059 \$16 \$12152 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14060 \$16 \$10348 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14062 \$16 \$10603 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14063 \$153 \$12019 \$10603 \$12130 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$14064 \$16 \$12236 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14065 \$16 \$10730 \$12012 \$12228 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$14066 \$153 \$12251 \$10634 \$12228 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$14067 \$153 \$12131 \$12019 \$12093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14069 \$153 \$11811 \$12251 \$12003 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14070 \$16 \$12003 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14071 \$16 \$12093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14072 \$16 \$10634 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14073 \$16 \$11898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14074 \$153 \$12132 \$12041 \$12003 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14075 \$153 \$12131 \$12229 \$12020 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14076 \$16 \$12003 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14077 \$16 \$12093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14079 \$16 \$12003 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14082 \$153 \$12063 \$12229 \$12252 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14083 \$16 \$12095 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14084 \$153 \$12092 \$12353 \$12252 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14085 \$153 \$12132 \$11810 \$12252 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14087 \$153 \$12185 \$12041 \$12158 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14088 \$16 \$12294 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14089 \$16 \$12236 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14090 \$16 \$12093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14093 \$153 \$12185 \$12057 \$12252 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14094 \$16 \$10744 \$12012 \$12023 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$14095 \$153 \$12186 \$11989 \$12093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14097 \$153 \$12253 \$11989 \$12152 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14098 \$16 \$12093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14099 \$16 \$12003 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14100 \$153 \$12186 \$12229 \$12094 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14102 \$16 \$10890 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14104 \$153 \$12187 \$11989 \$12095 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14105 \$16 \$12152 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14106 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$14107 \$153 \$12187 \$12353 \$12094 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14108 \$16 \$12158 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14109 \$16 \$12095 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14111 \$16 \$12230 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14112 \$16 \$10744 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14114 \$153 \$12171 \$12014 \$12158 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14116 \$153 \$12254 \$12014 \$12236 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14117 \$153 \$12171 \$12057 \$12004 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14118 \$153 \$12273 \$12208 \$12004 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14120 \$16 \$10555 \$16 \$153 \$12004 VNB sky130_fd_sc_hd__inv_1
X$14121 \$16 \$12158 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14123 \$16 \$12236 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14124 \$153 \$12188 \$12014 \$12093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14125 \$16 \$10555 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14126 \$153 \$12188 \$12229 \$12004 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14127 \$153 \$12207 \$12096 \$12093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14128 \$16 \$10413 \$12015 \$12133 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$14129 \$153 \$12153 \$12096 \$12095 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14131 \$16 \$12093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14133 \$153 \$12207 \$12229 \$12005 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14134 \$153 \$12153 \$12353 \$12005 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14135 \$153 \$12255 \$12208 \$12005 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14137 \$153 \$12097 \$11810 \$12005 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14139 \$153 \$12237 \$12209 \$12005 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14141 \$16 \$10413 \$16 \$153 \$12005 VNB sky130_fd_sc_hd__inv_1
X$14142 \$16 \$10413 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14143 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$14145 \$153 \$12098 \$12172 \$12095 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14146 \$153 \$12210 \$12172 \$12093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14147 \$16 \$12093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14148 \$16 \$12095 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14149 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$14150 \$16 \$10621 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14151 \$16 \$10621 \$16 \$153 \$12006 VNB sky130_fd_sc_hd__inv_1
X$14153 \$153 \$12211 \$12172 \$12003 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14154 \$153 \$12189 \$12172 \$12158 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14155 \$153 \$12211 \$11810 \$12006 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14156 \$153 \$12189 \$12057 \$12006 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14157 \$16 \$12158 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14160 \$16 \$12003 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14161 \$153 \$8364 \$12003 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$14162 \$16 \$10682 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14164 \$16 \$10732 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14165 \$16 \$11994 \$10667 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$14166 \$16 \$11994 \$10624 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$14167 \$16 \$11994 \$10706 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$14168 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$14169 \$16 \$8364 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14170 \$16 \$12016 \$11888 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$14171 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$14172 \$16 \$12016 \$11720 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$14173 \$153 \$9747 \$12095 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$14174 \$16 \$10730 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14176 \$153 \$9138 \$12093 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$14177 \$16 \$11805 \$12190 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$14178 \$16 \$9747 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14179 \$153 \$10179 \$8340 \$12208 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14180 \$16 \$9138 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14182 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14184 \$153 \$10151 \$8340 \$12134 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14186 \$16 \$12295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14187 \$153 \$12212 \$12191 \$12295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14188 \$153 \$12191 \$10603 \$12082 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$14191 \$153 \$12256 \$12191 \$12259 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14192 \$16 \$10348 \$16 \$153 \$12135 VNB sky130_fd_sc_hd__inv_1
X$14193 \$16 \$12296 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14194 \$153 \$12100 \$12068 \$12135 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14195 \$16 \$10348 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14196 \$16 \$12259 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14198 \$153 \$12173 \$12363 \$12154 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14199 \$153 \$12257 \$12191 \$12160 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14202 \$16 \$12083 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14203 \$153 \$12102 \$12174 \$12135 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14204 \$153 \$12257 \$12028 \$12135 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14205 \$16 \$10539 \$12159 \$12026 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$14206 \$16 \$12160 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14208 \$16 \$11757 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14209 \$153 \$12136 \$11996 \$12160 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14210 \$153 \$12136 \$12028 \$12238 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14213 \$16 \$10539 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14214 \$153 \$12239 \$12307 \$12238 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14215 \$16 \$10539 \$16 \$153 \$12238 VNB sky130_fd_sc_hd__inv_1
X$14216 \$16 \$12160 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14218 \$153 \$12137 \$11996 \$12083 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14219 \$153 \$12213 \$11996 \$12101 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14221 \$153 \$12137 \$12174 \$12238 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14222 \$153 \$12213 \$12476 \$12238 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14223 \$16 \$12083 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14224 \$16 \$12101 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14225 \$153 \$12105 \$12070 \$12160 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14226 \$153 \$12258 \$12070 \$12101 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14227 \$16 \$12160 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14229 \$153 \$12214 \$12070 \$12241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14230 \$16 \$12101 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14231 \$16 \$10890 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14232 \$153 \$12192 \$12070 \$12044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14233 \$16 \$12044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14234 \$153 \$12106 \$12174 \$12104 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14235 \$16 \$12083 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14236 \$16 \$10555 \$12161 \$12138 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$14238 \$153 \$12192 \$12068 \$12104 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14240 \$153 \$12193 \$12084 \$12083 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14241 \$153 \$12231 \$12155 \$12104 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14243 \$153 \$12045 \$10686 \$11660 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14244 \$153 \$12194 \$12084 \$12044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14245 \$16 \$10555 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14247 \$153 \$12193 \$12174 \$12071 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14248 \$153 \$12139 \$12084 \$12101 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14249 \$153 \$12194 \$12068 \$12071 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14250 \$153 \$12107 \$12028 \$12071 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14251 \$16 \$12044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14253 \$16 \$10621 \$16 \$153 \$12007 VNB sky130_fd_sc_hd__inv_1
X$14256 \$153 \$12215 \$12085 \$12295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14257 \$153 \$12139 \$12476 \$12071 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14258 \$16 \$12101 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14259 \$16 \$10621 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14260 \$16 \$12295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14261 \$153 \$12029 \$12085 \$12044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14262 \$153 \$12215 \$12155 \$12007 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14264 \$16 \$12044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14266 \$16 \$12259 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14267 \$153 \$12108 \$12174 \$12007 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14269 \$153 \$12308 \$10682 \$12260 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$14270 \$153 \$12030 \$12086 \$12101 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14271 \$16 \$10682 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14272 \$16 \$11488 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14274 \$153 \$12240 \$12359 \$11869 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14276 \$16 \$12101 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14278 \$16 \$10605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14279 \$16 \$10413 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14280 \$16 \$12083 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14281 \$16 \$11814 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14283 \$153 \$12261 \$12086 \$12241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14284 \$153 \$12195 \$12086 \$12160 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14285 \$153 \$12109 \$12068 \$11869 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14286 \$16 \$12241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14287 \$16 \$11164 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14289 \$153 \$12195 \$12028 \$11869 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14290 \$16 \$12160 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14291 \$153 \$8320 \$12259 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$14292 \$16 \$12190 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14293 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$14294 \$16 \$11814 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14295 \$153 \$12242 \$12068 \$12378 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14296 \$153 \$10383 \$12295 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$14299 \$16 \$8320 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14300 \$153 \$12072 \$11806 \$10605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14301 \$153 \$9747 \$12115 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$14302 \$153 \$11970 \$10344 \$11906 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14305 \$153 \$8364 \$12326 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$14306 \$153 \$8863 \$8340 \$12155 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14307 \$153 \$8523 \$8340 \$12363 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14308 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14310 \$153 \$10262 \$8340 \$12309 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14311 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14312 \$153 \$9885 \$8340 \$12582 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14313 \$153 \$11768 \$10417 \$11724 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14314 \$16 \$8568 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14315 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14318 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14319 \$153 \$10181 \$8340 \$12264 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14320 \$153 \$10253 \$8340 \$12603 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14322 \$153 \$11603 \$10417 \$11207 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14323 \$153 \$153 \$12217 \$12243 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14324 \$153 \$153 \$12110 \$12243 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14327 \$153 \$153 \$12165 \$12243 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14328 \$16 \$16 \$153 VNB sky130_fd_sc_hd__conb_1
X$14329 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14331 \$153 \$8539 \$8340 \$12359 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14332 \$153 \$8619 \$8340 \$12307 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14334 \$153 \$12196 \$12175 \$12219 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14337 \$153 \$12196 \$12110 \$12216 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14338 \$153 \$12262 \$12175 \$12115 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14339 \$153 \$11700 \$10472 \$11513 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14340 \$16 \$12162 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14341 \$16 \$12164 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14342 \$16 \$11930 \$11378 \$12008 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$14344 \$153 \$12197 \$12175 \$12164 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14345 \$16 \$10739 \$16 \$153 \$12216 VNB sky130_fd_sc_hd__inv_1
X$14346 \$153 \$11843 \$10833 \$11513 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14347 \$153 \$12197 \$12217 \$12216 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14348 \$153 \$11742 \$12198 \$12048 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$14349 \$16 \$12032 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14350 \$16 \$12009 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14352 \$153 \$12244 \$12603 \$12216 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14353 \$16 \$10578 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14354 \$16 \$12198 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14355 \$16 \$11013 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14357 \$16 \$12164 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14358 \$16 \$12219 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14359 \$153 \$12199 \$12163 \$12164 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14360 \$153 \$12263 \$12163 \$12219 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14365 \$153 \$12199 \$12217 \$12156 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14366 \$153 \$11880 \$12169 \$12112 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$14367 \$16 \$12297 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14368 \$153 \$12218 \$12163 \$12115 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14369 \$153 \$12281 \$12165 \$12156 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14370 \$16 \$12115 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14371 \$16 \$10736 \$16 \$153 \$12156 VNB sky130_fd_sc_hd__inv_1
X$14374 \$153 \$12218 \$12234 \$12156 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14375 \$153 \$12163 \$12220 \$12176 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$14376 \$16 \$12233 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14377 \$16 \$12169 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14379 \$16 \$10736 \$12166 \$12176 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$14380 \$16 \$12220 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14382 \$16 \$12219 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14383 \$16 \$10661 \$12166 \$12140 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$14384 \$153 \$12114 \$12113 \$12219 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14385 \$16 \$10661 \$16 \$153 \$12200 VNB sky130_fd_sc_hd__inv_1
X$14387 \$153 \$12201 \$12113 \$12115 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14388 \$153 \$12201 \$12234 \$12200 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14389 \$153 \$12202 \$12075 \$12115 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14390 \$153 \$12282 \$12264 \$12200 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14392 \$16 \$12233 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14395 \$153 \$12202 \$12234 \$11999 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14396 \$153 \$12141 \$12075 \$12219 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14397 \$153 \$12283 \$12217 \$11999 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14398 \$16 \$10649 \$12166 \$12116 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$14399 \$16 \$10597 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14400 \$16 \$12219 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14401 \$153 \$12221 \$12177 \$12219 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14403 \$16 \$12115 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14405 \$153 \$12203 \$12177 \$12115 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14406 \$153 \$12203 \$12234 \$12117 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14408 \$153 \$12204 \$10852 \$12222 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$14409 \$16 \$10853 \$12166 \$12222 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$14411 \$16 \$12298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14414 \$153 \$12265 \$12118 \$12298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14416 \$153 \$12142 \$12118 \$12219 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14417 \$153 \$12142 \$12110 \$12246 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14418 \$16 \$10852 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14419 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$14420 \$16 \$10529 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14421 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$14423 \$16 \$10529 \$12166 \$12205 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$14424 \$16 \$12164 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14425 \$16 \$12115 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14427 \$153 \$12206 \$12118 \$12115 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14428 \$153 \$12223 \$12118 \$12164 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14429 \$153 \$12206 \$12234 \$12246 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14430 \$16 \$10409 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14431 \$16 \$10853 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14432 \$16 \$10383 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14434 \$153 \$12223 \$12217 \$12246 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14435 \$16 \$12167 \$10960 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$14436 \$16 \$12167 \$10852 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$14437 \$16 \$12167 \$12050 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$14438 \$16 \$8320 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14439 \$16 \$12167 \$10860 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$14440 \$16 \$12167 \$12245 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$14441 \$16 \$12167 \$12220 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$14442 \$153 \$8320 \$12299 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$14444 \$16 \$12168 \$16 \$153 \$12167 VNB sky130_fd_sc_hd__clkbuf_2
X$14445 \$16 \$12167 \$10981 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$14446 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14448 \$153 \$8416 \$12010 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$14449 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14450 \$153 \$8808 \$8340 \$12339 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14451 \$16 \$8416 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14452 \$16 \$12119 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14453 \$16 \$11148 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14454 \$16 \$12339 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14455 \$16 \$10311 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14456 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14457 \$153 \$10311 \$12384 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$14459 \$153 \$7995 \$8340 \$12227 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14461 \$153 \$12224 \$12178 \$11983 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14462 \$16 \$11983 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14463 \$16 \$12227 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14464 \$16 \$12287 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14465 \$16 \$12010 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14468 \$153 \$12143 \$12178 \$12010 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14469 \$153 \$12224 \$11881 \$12247 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14470 \$153 \$12248 \$12339 \$12247 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14471 \$153 \$12143 \$11942 \$12247 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14473 \$16 \$12384 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14474 \$153 \$12144 \$12178 \$12384 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14475 \$16 \$12120 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14477 \$153 \$12225 \$12178 \$12120 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14478 \$153 \$12144 \$12179 \$12247 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14479 \$153 \$12225 \$12182 \$12247 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14481 \$16 \$11983 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14482 \$16 \$12010 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14483 \$153 \$12122 \$12170 \$11983 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14485 \$153 \$12145 \$12170 \$12010 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14486 \$153 \$12249 \$12371 \$12121 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14487 \$153 \$12123 \$12170 \$12120 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14488 \$16 \$12384 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14489 \$16 \$10739 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14490 \$16 \$12351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14492 \$153 \$12266 \$12170 \$12351 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14493 \$16 \$10739 \$16 \$153 \$12121 VNB sky130_fd_sc_hd__inv_1
X$14494 \$16 \$12198 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14496 \$153 \$11681 \$12169 \$12053 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$14497 \$16 \$12169 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14499 \$16 \$10649 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14500 \$16 \$12351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14502 \$153 \$12226 \$12087 \$12351 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14503 \$16 \$12299 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14505 \$153 \$12035 \$12087 \$12299 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14506 \$153 \$12266 \$12119 \$12121 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14507 \$153 \$12180 \$12220 \$12146 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$14508 \$16 \$10649 \$12018 \$12125 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$14509 \$16 \$12303 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14513 \$16 \$11983 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14514 \$153 \$12349 \$12179 \$12147 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14515 \$153 \$12054 \$12087 \$11983 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14516 \$16 \$10736 \$16 \$153 \$12302 VNB sky130_fd_sc_hd__inv_1
X$14518 \$16 \$12010 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14519 \$153 \$12267 \$12180 \$12010 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14520 \$16 \$10649 \$16 \$153 \$12147 VNB sky130_fd_sc_hd__inv_1
X$14521 \$16 \$10661 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14522 \$16 \$10649 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14525 \$153 \$12055 \$10815 \$11730 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14526 \$153 \$12268 \$12180 \$11983 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14528 \$16 \$12299 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14529 \$153 \$12157 \$12088 \$12299 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14530 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$14531 \$16 \$10661 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14535 \$153 \$12157 \$12371 \$12127 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14536 \$16 \$12120 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14537 \$153 \$12290 \$12179 \$12127 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14538 \$16 \$10661 \$16 \$153 \$12127 VNB sky130_fd_sc_hd__inv_1
X$14541 \$153 \$12089 \$10852 \$12128 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$14542 \$16 \$10597 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14543 \$16 \$12299 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14544 \$153 \$12181 \$12089 \$12299 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14546 \$16 \$10852 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14548 \$153 \$12181 \$12371 \$11958 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14549 \$153 \$12269 \$12089 \$12384 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14550 \$16 \$12384 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14551 \$153 \$12148 \$12089 \$12120 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14552 \$16 \$12303 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14553 \$16 \$10853 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14555 \$16 \$10960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14558 \$153 \$12148 \$12182 \$11958 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14559 \$16 \$12287 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14560 \$153 \$12292 \$12227 \$11958 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14562 \$16 \$12120 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14564 \$16 \$10529 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14565 \$153 \$12270 \$12037 \$12120 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14566 \$16 \$11798 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14568 \$153 \$12129 \$11881 \$12011 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14570 \$153 \$12270 \$12182 \$12011 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14571 \$153 \$12271 \$12037 \$12287 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14573 \$16 \$12299 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14574 \$153 \$12149 \$12037 \$12299 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14575 \$16 \$12351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14576 \$153 \$12235 \$12119 \$12011 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14578 \$153 \$12235 \$12037 \$12351 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14579 \$153 \$12149 \$12371 \$12011 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14580 \$153 \$11386 \$10466 \$11390 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14581 \$153 \$11927 \$10642 \$11926 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14582 \$153 \$11320 \$10815 \$11390 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14583 \$153 \$11714 \$10694 \$11926 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14585 \$16 \$11390 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14586 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$14587 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$14588 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$14589 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$14590 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$14591 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$14592 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$14594 \$153 \$1728 \$1465 \$263 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14595 \$153 \$1785 \$1547 \$1762 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14596 \$153 \$1786 \$1792 \$1762 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14597 \$153 \$1629 \$102 \$1535 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14599 \$153 \$1728 \$234 \$1535 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14600 \$16 \$710 \$1430 \$1729 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$14602 \$16 \$1430 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14603 \$153 \$1683 \$1465 \$249 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14604 \$16 \$264 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14605 \$153 \$2193 \$753 \$1729 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$14608 \$16 \$264 \$1430 \$1814 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$14609 \$153 \$1683 \$377 \$1535 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14611 \$153 \$1546 \$1774 \$1658 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14612 \$153 \$1684 \$2009 \$1669 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14613 \$16 \$1658 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14614 \$153 \$1257 \$1595 \$1685 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$14615 \$16 \$1480 \$1168 \$1685 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$14618 \$153 \$1787 \$1943 \$1537 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14619 \$153 \$1656 \$1257 \$263 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14620 \$153 \$1788 \$2252 \$1537 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14621 \$153 \$1790 \$1547 \$1789 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14623 \$16 \$754 \$1430 \$1730 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$14624 \$153 \$1763 \$662 \$1730 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$14626 \$153 \$1656 \$234 \$1106 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14628 \$153 \$1326 \$1686 \$1498 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$14629 \$153 \$1791 \$1792 \$1537 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14631 \$16 \$582 \$1522 \$1764 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$14632 \$153 \$1548 \$1326 \$184 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14634 \$16 \$1687 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14635 \$153 \$1774 \$430 \$1764 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$14636 \$153 \$1657 \$30 \$1327 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14637 \$153 \$1888 \$541 \$1731 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$14638 \$16 \$279 \$1522 \$1731 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$14639 \$16 \$184 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14641 \$153 \$1550 \$1249 \$184 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14643 \$16 \$58 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14644 \$153 \$1794 \$1792 \$1793 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14645 \$153 \$1963 \$454 \$1765 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$14646 \$153 \$1630 \$30 \$1250 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14647 \$153 \$1258 \$1553 \$1570 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$14649 \$16 \$280 \$1430 \$1765 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$14651 \$16 \$1553 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14652 \$153 \$1766 \$1525 \$1732 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$14653 \$16 \$323 \$1430 \$1732 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$14655 \$16 \$58 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14656 \$153 \$1452 \$394 \$1454 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14657 \$16 \$1795 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14658 \$153 \$1747 \$1766 \$1687 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14660 \$153 \$1500 \$234 \$1191 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14662 \$153 \$1434 \$561 \$1454 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14663 \$153 \$1747 \$1792 \$1767 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14664 \$153 \$1733 \$1675 \$1658 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14665 \$16 \$323 \$16 \$153 \$1767 VNB sky130_fd_sc_hd__inv_1
X$14666 \$16 \$1687 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14667 \$16 \$58 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14669 \$16 \$1795 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14671 \$16 \$1687 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14672 \$153 \$1840 \$1792 \$1796 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14673 \$16 \$1658 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14674 \$16 \$1348 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14675 \$16 \$1525 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14676 \$153 \$1675 \$535 \$1688 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$14677 \$16 \$356 \$1430 \$1688 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$14679 \$153 \$1676 \$684 \$1734 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$14682 \$16 \$380 \$1522 \$1734 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$14683 \$16 \$1687 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14684 \$153 \$1748 \$1676 \$1687 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14685 \$153 \$1689 \$1676 \$1658 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14686 \$16 \$380 \$16 \$153 \$1670 VNB sky130_fd_sc_hd__inv_1
X$14687 \$153 \$1689 \$1547 \$1670 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14688 \$16 \$356 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14691 \$16 \$684 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14692 \$16 \$1687 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14693 \$16 \$1658 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14694 \$153 \$1749 \$1797 \$1687 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14695 \$16 \$380 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14696 \$16 \$1522 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14697 \$16 \$58 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14698 \$16 \$351 \$1522 \$1690 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$14699 \$153 \$1691 \$1815 \$1671 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14700 \$153 \$1797 \$505 \$1690 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$14701 \$16 \$184 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14703 \$16 \$1552 \$1047 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$14704 \$16 \$1552 \$535 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$14705 \$16 \$1552 \$753 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$14707 \$153 \$1775 \$184 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$14708 \$16 \$1552 \$662 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$14709 \$16 \$1331 \$1659 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$14710 \$16 \$1625 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14711 \$16 \$505 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14713 \$16 \$1626 \$1686 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$14714 \$16 \$1626 \$1503 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$14715 \$16 \$1626 \$1208 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$14719 \$16 \$1626 \$1576 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$14720 \$16 \$1776 \$16 \$153 \$280 VNB sky130_fd_sc_hd__clkbuf_2
X$14721 \$16 \$349 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14722 \$16 \$1798 \$16 \$153 \$323 VNB sky130_fd_sc_hd__clkbuf_2
X$14723 \$153 \$1918 \$58 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$14724 \$16 \$1777 \$1799 \$1816 \$1768 \$16 \$153 \$1778 VNB
+ sky130_fd_sc_hd__and4_2
X$14725 \$16 \$1800 \$16 \$153 \$356 VNB sky130_fd_sc_hd__clkbuf_2
X$14726 \$16 \$1778 \$16 \$153 \$754 VNB sky130_fd_sc_hd__clkbuf_2
X$14727 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14729 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14731 \$153 \$1750 \$1482 \$377 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14733 \$153 \$1735 \$1482 \$349 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14734 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14735 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14736 \$16 \$1801 \$16 \$153 \$351 VNB sky130_fd_sc_hd__clkbuf_2
X$14737 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14738 \$153 \$1692 \$1482 \$30 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14740 \$16 \$280 \$1292 \$1817 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$14742 \$153 \$1802 \$1482 \$102 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14743 \$16 \$102 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14744 \$16 \$30 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14745 \$16 \$1480 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14746 \$16 \$1480 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14747 \$153 \$1632 \$35 \$1633 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14748 \$153 \$1693 \$54 \$1633 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14749 \$153 \$1751 \$1482 \$59 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14750 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14752 \$16 \$280 \$16 \$153 \$1864 VNB sky130_fd_sc_hd__inv_1
X$14753 \$16 \$264 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14754 \$16 \$454 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14755 \$153 \$1634 \$346 \$1633 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14756 \$153 \$1505 \$253 \$1633 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14757 \$16 \$280 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14758 \$153 \$1694 \$1919 \$1845 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14759 \$16 \$1923 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14760 \$16 \$662 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14761 \$16 \$1292 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14764 \$153 \$1779 \$662 \$1736 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$14765 \$16 \$754 \$1292 \$1736 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$14767 \$153 \$1575 \$104 \$1633 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14768 \$153 \$1804 \$1779 \$1923 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14769 \$16 \$1348 \$979 \$1636 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$14770 \$16 \$1348 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14772 \$153 \$1695 \$1779 \$1805 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14773 \$153 \$1694 \$1471 \$1864 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14774 \$153 \$1695 \$1703 \$1483 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14775 \$153 \$1803 \$1924 \$1483 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14776 \$16 \$1805 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14779 \$153 \$1769 \$1806 \$1483 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14780 \$16 \$1404 \$979 \$1662 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$14781 \$153 \$1697 \$753 \$1696 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$14782 \$153 \$1804 \$1895 \$1483 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14784 \$16 \$1923 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14785 \$16 \$710 \$1292 \$1696 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$14786 \$153 \$1818 \$1697 \$1805 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14787 \$16 \$979 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14789 \$153 \$1637 \$1334 \$212 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14790 \$16 \$1805 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14792 \$153 \$1819 \$1697 \$1845 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14793 \$153 \$1698 \$1895 \$1866 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14794 \$16 \$212 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14797 \$16 \$1328 \$979 \$1663 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$14798 \$153 \$1820 \$1525 \$1638 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$14799 \$153 \$1843 \$1471 \$1844 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14800 \$153 \$1700 \$535 \$1699 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$14802 \$16 \$356 \$1292 \$1699 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$14803 \$153 \$1821 \$1820 \$1805 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14805 \$16 \$979 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14806 \$153 \$1577 \$35 \$1335 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14808 \$153 \$1807 \$1700 \$1923 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14809 \$153 \$1701 \$1421 \$212 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14810 \$16 \$356 \$16 \$153 \$1822 VNB sky130_fd_sc_hd__inv_1
X$14811 \$153 \$1701 \$347 \$1335 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14813 \$153 \$1639 \$1700 \$1845 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14814 \$16 \$212 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14815 \$16 \$1328 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14816 \$153 \$1672 \$1472 \$212 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14817 \$153 \$1770 \$684 \$1823 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$14819 \$153 \$1702 \$1703 \$1822 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14821 \$16 \$380 \$16 \$153 \$1752 VNB sky130_fd_sc_hd__inv_1
X$14822 \$153 \$1753 \$1770 \$1923 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14823 \$153 \$1672 \$347 \$1410 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14824 \$16 \$212 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14826 \$16 \$1923 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14827 \$16 \$351 \$1966 \$1824 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$14828 \$153 \$1641 \$1472 \$293 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14831 \$153 \$1754 \$1770 \$1805 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14832 \$153 \$1846 \$1471 \$1752 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14833 \$153 \$1825 \$1780 \$1923 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14834 \$16 \$351 \$16 \$153 \$1704 VNB sky130_fd_sc_hd__inv_1
X$14835 \$16 \$293 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14836 \$16 \$1805 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14840 \$153 \$1673 \$293 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$14842 \$153 \$1755 \$1780 \$1845 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14843 \$16 \$1965 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14844 \$16 \$1673 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14845 \$16 \$1923 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14847 \$153 \$153 \$347 \$1487 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14848 \$16 \$1845 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14851 \$153 \$1825 \$1895 \$1704 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14853 \$153 \$1677 \$209 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$14855 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14856 \$153 \$1737 \$1482 \$35 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14857 \$16 \$1677 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14859 \$16 \$1775 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14860 \$153 \$1678 \$212 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$14861 \$153 \$1775 \$241 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$14862 \$153 \$1918 \$424 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$14863 \$16 \$1678 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14864 \$16 \$1918 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14865 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14867 \$153 \$1826 \$1482 \$253 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14868 \$153 \$1705 \$1482 \$215 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14869 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14870 \$16 \$215 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14872 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14873 \$153 \$1848 \$1712 \$1540 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14875 \$153 \$1706 \$1482 \$346 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14876 \$153 \$2407 \$1482 \$266 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14877 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14878 \$16 \$1756 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14879 \$16 \$1969 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14881 \$153 \$1644 \$1781 \$1969 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14882 \$153 \$1559 \$1183 \$241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14883 \$153 \$1808 \$1712 \$1679 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14884 \$16 \$241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14886 \$16 \$1543 \$1446 \$1739 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$14888 \$153 \$1183 \$1760 \$1739 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$14891 \$16 \$399 \$1929 \$1740 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$14892 \$153 \$1741 \$1268 \$424 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14893 \$153 \$1268 \$1628 \$1512 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$14895 \$16 \$1566 \$16 \$153 \$1396 VNB sky130_fd_sc_hd__inv_1
X$14896 \$16 \$1756 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14897 \$153 \$1338 \$1933 \$1580 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$14899 \$153 \$1741 \$353 \$1396 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14900 \$153 \$1850 \$1712 \$1771 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14901 \$153 \$1616 \$1338 \$241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14902 \$153 \$1827 \$1338 \$424 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14904 \$16 \$1585 \$16 \$153 \$1811 VNB sky130_fd_sc_hd__inv_1
X$14905 \$153 \$1680 \$353 \$1456 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14907 \$153 \$1809 \$1558 \$1771 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14908 \$153 \$1253 \$1708 \$1707 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$14909 \$153 \$1828 \$1613 \$1771 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14911 \$153 \$1560 \$1253 \$424 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14912 \$16 \$241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14914 \$153 \$1645 \$1253 \$241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14915 \$153 \$1709 \$1712 \$1674 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14916 \$16 \$1518 \$16 \$153 \$1541 VNB sky130_fd_sc_hd__inv_1
X$14918 \$153 \$1270 \$1647 \$1742 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$14919 \$16 \$1518 \$1446 \$1707 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$14921 \$16 \$1514 \$1446 \$1742 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$14923 \$153 \$1757 \$1270 \$241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14924 \$153 \$1680 \$1270 \$424 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14925 \$16 \$1514 \$16 \$153 \$1456 VNB sky130_fd_sc_hd__inv_1
X$14926 \$16 \$241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14927 \$16 \$591 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14928 \$16 \$1446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14929 \$16 \$1758 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14930 \$16 \$1708 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14932 \$153 \$1710 \$1868 \$1542 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14933 \$153 \$1810 \$1613 \$1674 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14935 \$153 \$1711 \$2438 \$1542 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14936 \$16 \$1758 \$1446 \$1829 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$14938 \$153 \$1648 \$1254 \$424 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14939 \$153 \$1713 \$1712 \$1542 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14941 \$153 \$1714 \$1715 \$1542 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14942 \$153 \$1903 \$608 \$1830 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$14943 \$16 \$1758 \$16 \$153 \$1412 VNB sky130_fd_sc_hd__inv_1
X$14945 \$16 \$424 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14946 \$153 \$1716 \$1320 \$424 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14947 \$153 \$1772 \$1613 \$1542 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14951 \$16 \$306 \$16 \$153 \$1759 VNB sky130_fd_sc_hd__inv_1
X$14952 \$16 \$608 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14953 \$153 \$1852 \$1558 \$1759 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14954 \$153 \$1320 \$1649 \$1717 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$14955 \$153 \$1757 \$388 \$1456 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14956 \$153 \$1646 \$266 \$1456 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14957 \$153 \$1239 \$112 \$1456 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14959 \$153 \$1424 \$1593 \$1584 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$14960 \$153 \$1616 \$388 \$1811 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14961 \$153 \$1455 \$266 \$1811 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14962 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14963 \$153 \$2166 \$1482 \$57 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14964 \$16 \$1879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14965 \$16 \$241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14966 \$16 \$724 \$16 \$153 \$1996 VNB sky130_fd_sc_hd__inv_1
X$14969 \$153 \$1681 \$1424 \$241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14970 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14971 \$16 \$1475 \$16 \$153 \$1229 VNB sky130_fd_sc_hd__inv_1
X$14972 \$153 \$1718 \$1482 \$23 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14973 \$153 \$1782 \$1831 \$1682 \$1970 \$1812 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$14975 \$16 \$1678 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14978 \$16 \$1677 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$14979 \$153 \$1681 \$388 \$1229 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$14980 \$153 \$1677 \$178 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$14981 \$16 \$1682 \$16 \$153 \$151 VNB sky130_fd_sc_hd__clkbuf_2
X$14982 \$153 \$1678 \$446 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$14984 \$16 \$1783 \$1459 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$14985 \$16 \$1783 \$1489 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$14988 \$16 \$1783 \$387 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$14990 \$153 \$1720 \$1482 \$398 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$14991 \$16 \$1783 \$631 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$14992 \$16 \$1783 \$558 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$14994 \$16 \$1721 \$16 \$153 \$1783 VNB sky130_fd_sc_hd__clkbuf_2
X$14995 \$16 \$1783 \$884 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$14997 \$16 \$1721 \$16 \$153 \$1832 VNB sky130_fd_sc_hd__clkbuf_2
X$14998 \$16 \$1482 \$16 \$153 \$1721 VNB sky130_fd_sc_hd__clkbuf_2
X$14999 \$16 \$1783 \$674 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$15000 \$16 \$1783 \$856 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$15001 \$16 \$1784 \$591 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$15003 \$16 \$1721 \$16 \$153 \$1784 VNB sky130_fd_sc_hd__clkbuf_2
X$15004 \$16 \$1784 \$595 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$15005 \$16 \$1564 \$1719 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$15006 \$16 \$1784 \$948 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$15007 \$16 \$1564 \$895 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$15008 \$16 \$1784 \$423 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$15009 \$16 \$1832 \$1627 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$15010 \$16 \$1784 \$1245 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$15011 \$16 \$63 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15012 \$16 \$1784 \$608 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$15013 \$153 \$1340 \$1760 \$1722 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$15014 \$16 \$1832 \$1708 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$15015 \$16 \$1832 \$1593 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$15016 \$16 \$1972 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15018 \$16 \$1860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15021 \$16 \$1543 \$1601 \$1722 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$15022 \$16 \$1585 \$1601 \$1773 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$15024 \$153 \$1565 \$1933 \$1773 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$15025 \$153 \$1587 \$23 \$1341 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15026 \$153 \$1618 \$371 \$1341 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15027 \$153 \$1620 \$1565 \$446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15028 \$16 \$1585 \$16 \$153 \$1651 VNB sky130_fd_sc_hd__inv_1
X$15030 \$153 \$1743 \$1565 \$178 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15032 \$153 \$1743 \$549 \$1651 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15034 \$153 \$1857 \$1565 \$509 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15036 \$153 \$1745 \$371 \$1491 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15039 \$153 \$1622 \$1628 \$1744 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$15040 \$16 \$1566 \$1601 \$1744 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$15041 \$153 \$1745 \$1622 \$509 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15042 \$153 \$1462 \$703 \$1491 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15043 \$153 \$1517 \$223 \$1491 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15044 \$16 \$178 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15046 \$16 \$1566 \$16 \$153 \$1491 VNB sky130_fd_sc_hd__inv_1
X$15047 \$153 \$1723 \$1622 \$178 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15048 \$16 \$446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15049 \$153 \$1652 \$1622 \$446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15050 \$153 \$1723 \$549 \$1491 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15051 \$16 \$1518 \$1601 \$1833 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$15052 \$16 \$1601 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15054 \$16 \$151 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15056 \$16 \$1601 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15057 \$16 \$591 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15058 \$16 \$446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15059 \$16 \$178 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15060 \$153 \$1653 \$1342 \$446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15061 \$153 \$1666 \$1342 \$178 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15062 \$16 \$1885 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15063 \$16 \$1518 \$16 \$153 \$1255 VNB sky130_fd_sc_hd__inv_1
X$15064 \$16 \$509 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15065 \$16 \$306 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15066 \$153 \$1302 \$1647 \$1859 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$15068 \$153 \$1666 \$549 \$1255 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15070 \$16 \$446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15071 \$153 \$1834 \$1302 \$509 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15072 \$153 \$1667 \$1302 \$446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15073 \$153 \$1667 \$393 \$1343 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15075 \$153 \$1592 \$703 \$1343 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15076 \$16 \$1514 \$16 \$153 \$1343 VNB sky130_fd_sc_hd__inv_1
X$15077 \$16 \$446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15078 \$153 \$1724 \$1492 \$446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15079 \$16 \$178 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15080 \$153 \$1725 \$1492 \$178 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15082 \$153 \$1725 \$549 \$1414 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15083 \$16 \$1599 \$16 \$153 \$1414 VNB sky130_fd_sc_hd__inv_1
X$15084 \$16 \$509 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15085 \$153 \$1623 \$1492 \$509 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15086 \$153 \$1724 \$393 \$1414 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15088 \$153 \$1568 \$1593 \$1655 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$15089 \$16 \$1758 \$1601 \$1835 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$15093 \$16 \$509 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15094 \$16 \$509 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15097 \$153 \$1746 \$1568 \$509 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15098 \$153 \$1668 \$1416 \$509 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15099 \$16 \$1475 \$16 \$153 \$1344 VNB sky130_fd_sc_hd__inv_1
X$15100 \$16 \$1758 \$16 \$153 \$1415 VNB sky130_fd_sc_hd__inv_1
X$15102 \$16 \$178 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15103 \$16 \$178 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15104 \$153 \$1761 \$1416 \$178 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15106 \$153 \$1726 \$1568 \$178 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15107 \$153 \$1761 \$549 \$1415 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15109 \$153 \$1727 \$1568 \$446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15110 \$16 \$446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15113 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$15114 \$153 \$1726 \$549 \$1344 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15115 \$153 \$1813 \$393 \$1415 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15116 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$15117 \$153 \$1727 \$393 \$1344 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15118 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$15119 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$15122 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$15124 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$15125 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$15126 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$15127 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$15130 \$153 \$11519 \$11499 \$10368 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15131 \$153 \$11286 \$11288 \$10368 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15132 \$16 \$10368 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15133 \$153 \$11362 \$10327 \$11232 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15134 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$15136 \$153 \$11418 \$11288 \$10200 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15137 \$153 \$11520 \$11499 \$10200 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15138 \$153 \$11419 \$11499 \$10367 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15139 \$153 \$11418 \$10088 \$11232 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15140 \$16 \$10646 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15142 \$16 \$10200 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15143 \$153 \$11288 \$11432 \$11363 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$15144 \$16 \$10367 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15145 \$16 \$10200 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15146 \$153 \$11465 \$11499 \$10476 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15147 \$153 \$11419 \$10330 \$11263 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15148 \$16 \$10476 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15149 \$16 \$11432 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15151 \$16 \$11289 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15154 \$153 \$11465 \$10705 \$11263 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15155 \$153 \$11420 \$11348 \$10200 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15157 \$16 \$10200 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15158 \$16 \$10427 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15159 \$153 \$11400 \$11348 \$10427 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15160 \$153 \$11420 \$10088 \$11265 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15163 \$153 \$11400 \$10327 \$11265 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15164 \$16 \$11369 \$11347 \$11523 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$15165 \$153 \$11466 \$11348 \$10295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15167 \$16 \$10367 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15168 \$153 \$11421 \$11348 \$10476 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15169 \$16 \$11369 \$16 \$153 \$11265 VNB sky130_fd_sc_hd__inv_1
X$15170 \$16 \$10295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15171 \$153 \$11421 \$10705 \$11265 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15173 \$153 \$11466 \$10276 \$11265 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15174 \$16 \$10476 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15176 \$153 \$11467 \$11271 \$10367 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15177 \$153 \$11422 \$11271 \$10476 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15178 \$153 \$11468 \$11271 \$10226 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15181 \$153 \$11467 \$10330 \$11191 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15182 \$16 \$10476 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15184 \$153 \$11424 \$11484 \$10200 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15185 \$153 \$11422 \$10705 \$11191 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15186 \$16 \$10226 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15187 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$15190 \$153 \$11524 \$11484 \$10368 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15191 \$153 \$11423 \$10327 \$11393 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15192 \$153 \$11424 \$10088 \$11393 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15193 \$16 \$10368 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15194 \$153 \$11525 \$11484 \$10646 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15195 \$16 \$11297 \$16 \$153 \$11191 VNB sky130_fd_sc_hd__inv_1
X$15196 \$16 \$11297 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15197 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$15199 \$16 \$11297 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15201 \$153 \$11401 \$10161 \$11393 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15202 \$153 \$11470 \$11484 \$10476 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15203 \$16 \$10646 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15204 \$153 \$11470 \$10705 \$11393 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15206 \$16 \$11485 \$11238 \$11486 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$15207 \$153 \$11365 \$10161 \$10954 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15209 \$153 \$11484 \$11637 \$11486 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$15210 \$16 \$11240 \$11238 \$11394 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$15211 \$153 \$11000 \$11856 \$11394 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$15212 \$153 \$11469 \$10276 \$11652 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15213 \$16 \$10200 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15214 \$16 \$11856 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15215 \$16 \$10427 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15217 \$153 \$11404 \$11425 \$10226 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15219 \$153 \$11426 \$11425 \$10427 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15220 \$153 \$11505 \$10330 \$11395 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15221 \$153 \$11426 \$10327 \$11395 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15222 \$16 \$10226 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15223 \$16 \$11637 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15224 \$153 \$11402 \$10705 \$11395 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15227 \$153 \$11403 \$11425 \$10646 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15228 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$15229 \$153 \$11403 \$10318 \$11395 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15230 \$16 \$10646 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15231 \$153 \$11404 \$10161 \$11395 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15232 \$153 \$11471 \$11425 \$10368 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15235 \$16 \$10974 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15236 \$16 \$11196 \$16 \$153 \$10825 VNB sky130_fd_sc_hd__clkbuf_2
X$15237 \$153 \$11471 \$10303 \$11395 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15238 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$15239 \$16 \$11350 \$16 \$153 \$10732 VNB sky130_fd_sc_hd__clkbuf_2
X$15240 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$15241 \$16 \$10368 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15242 \$16 \$11351 \$16 \$153 \$11427 VNB sky130_fd_sc_hd__clkbuf_2
X$15244 \$153 \$11527 \$11429 \$11427 \$11428 \$11430 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$15245 \$16 \$11244 \$16 \$153 \$11428 VNB sky130_fd_sc_hd__clkbuf_2
X$15246 \$16 \$11119 \$16 \$153 \$11429 VNB sky130_fd_sc_hd__clkbuf_2
X$15248 \$16 \$11111 \$16 \$153 \$11180 VNB sky130_fd_sc_hd__clkbuf_2
X$15249 \$153 \$11428 \$11429 \$11506 \$11430 \$11427 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$15250 \$16 \$11294 \$16 \$153 \$10621 VNB sky130_fd_sc_hd__clkbuf_2
X$15251 \$16 \$11352 \$16 \$153 \$10747 VNB sky130_fd_sc_hd__clkbuf_2
X$15252 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$15253 \$16 \$11111 \$16 \$153 \$11430 VNB sky130_fd_sc_hd__clkbuf_2
X$15254 \$16 \$11119 \$16 \$153 \$11507 VNB sky130_fd_sc_hd__clkbuf_2
X$15256 \$16 \$11272 \$11296 \$11273 \$153 \$11199 \$16 VNB
+ sky130_fd_sc_hd__and3b_4
X$15258 \$153 \$11528 \$11507 \$11529 \$11508 \$11561 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$15260 \$16 \$11244 \$16 \$153 \$11508 VNB sky130_fd_sc_hd__clkbuf_2
X$15262 \$16 \$11432 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15263 \$153 \$11120 \$11432 \$11405 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$15264 \$16 \$11289 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15265 \$16 \$11289 \$11275 \$11405 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$15267 \$153 \$11530 \$11500 \$10526 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15268 \$153 \$11433 \$11120 \$10605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15271 \$153 \$11487 \$11500 \$10338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15272 \$153 \$11433 \$10686 \$11200 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15273 \$153 \$11434 \$10686 \$11396 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15274 \$16 \$10526 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15275 \$16 \$10338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15276 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$15277 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$15278 \$153 \$11472 \$11500 \$10470 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15280 \$153 \$11367 \$10309 \$11200 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15281 \$153 \$11368 \$10247 \$11200 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15282 \$153 \$11472 \$10247 \$11396 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15283 \$16 \$10470 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15284 \$16 \$10470 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15285 \$153 \$11370 \$11121 \$10606 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15287 \$16 \$11369 \$11275 \$11532 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$15289 \$153 \$11473 \$11121 \$10605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15290 \$153 \$11473 \$10686 \$11112 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15292 \$153 \$11340 \$11121 \$10470 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15293 \$16 \$10606 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15294 \$16 \$10605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15295 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$15298 \$16 \$11369 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15300 \$16 \$11123 \$16 \$153 \$11275 VNB sky130_fd_sc_hd__clkbuf_2
X$15301 \$153 \$11533 \$11435 \$10298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15302 \$153 \$11436 \$11435 \$10605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15303 \$16 \$10298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15304 \$16 \$10605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15305 \$153 \$11437 \$11435 \$10606 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15306 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$15309 \$153 \$11509 \$10309 \$11397 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15310 \$153 \$11437 \$10344 \$11397 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15311 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$15312 \$153 \$11534 \$11435 \$10526 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15313 \$16 \$10606 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15314 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$15315 \$16 \$10526 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15317 \$153 \$11438 \$11435 \$10382 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15318 \$153 \$11474 \$11435 \$10514 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15319 \$16 \$10382 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15320 \$153 \$11438 \$10098 \$11397 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15322 \$153 \$11389 \$11439 \$10338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15323 \$16 \$10514 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15325 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$15326 \$153 \$11475 \$11439 \$10526 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15327 \$153 \$11389 \$10309 \$11398 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15328 \$153 \$11406 \$10247 \$11398 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15329 \$153 \$11475 \$10516 \$11398 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15330 \$16 \$10338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15333 \$16 \$10605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15334 \$16 \$10526 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15335 \$16 \$11194 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15337 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$15338 \$16 \$11488 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15339 \$16 \$11488 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15340 \$153 \$11440 \$11439 \$10382 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15341 \$153 \$11476 \$11439 \$10514 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15343 \$16 \$10514 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15344 \$153 \$11440 \$10098 \$11398 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15345 \$16 \$11164 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15347 \$153 \$11476 \$10538 \$11398 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15349 \$16 \$11240 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15350 \$153 \$11302 \$10098 \$11061 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15351 \$16 \$11240 \$11164 \$11535 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$15353 \$153 \$11441 \$11276 \$10526 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15354 \$16 \$11431 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15355 \$153 \$11407 \$10344 \$11205 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15357 \$16 \$10470 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15358 \$153 \$11441 \$10516 \$11205 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15359 \$16 \$10526 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15360 \$16 \$11164 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15361 \$16 \$11240 \$16 \$153 \$11205 VNB sky130_fd_sc_hd__inv_1
X$15362 \$153 \$11536 \$11276 \$10338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15363 \$153 \$11371 \$10401 \$11205 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15365 \$16 \$10605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15366 \$16 \$10382 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15367 \$153 \$11208 \$11431 \$11372 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$15368 \$16 \$10338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15370 \$153 \$11510 \$10538 \$11205 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15371 \$16 \$10514 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15373 \$153 \$11442 \$11208 \$10382 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15374 \$16 \$10382 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15375 \$16 \$10382 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15376 \$153 \$11477 \$11208 \$10606 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15379 \$153 \$11442 \$10098 \$11268 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15380 \$153 \$11477 \$10344 \$11268 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15381 \$16 \$11164 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15382 \$16 \$10606 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15383 \$16 \$10338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15384 \$153 \$11443 \$11208 \$10338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15385 \$16 \$11488 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15386 \$16 \$11488 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15388 \$153 \$11511 \$10309 \$11906 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15391 \$153 \$11443 \$10309 \$11268 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15392 \$153 \$11353 \$11208 \$10470 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15393 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$15394 \$16 \$10735 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15395 \$153 \$10828 \$11501 \$10735 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15397 \$153 \$11408 \$10471 \$11207 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15399 \$16 \$10300 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15400 \$16 \$10473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15401 \$153 \$11165 \$11501 \$10473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15402 \$16 \$11207 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15404 \$153 \$11128 \$11501 \$10578 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15405 \$16 \$10611 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15406 \$16 \$12234 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15407 \$16 \$12217 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15408 \$16 \$10578 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15410 \$16 \$11399 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15411 \$153 \$10976 \$11501 \$10386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15414 \$16 \$11374 \$11127 \$11538 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$15415 \$153 \$11489 \$10833 \$11065 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15416 \$16 \$10386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15417 \$153 \$11512 \$10417 \$11065 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15418 \$16 \$10578 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15419 \$153 \$11375 \$10501 \$11065 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15420 \$153 \$11489 \$11185 \$10611 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15422 \$153 \$11444 \$11185 \$10578 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15423 \$16 \$10551 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15424 \$16 \$10300 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15425 \$16 \$10611 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15427 \$153 \$11409 \$10471 \$11065 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15429 \$153 \$11490 \$10417 \$11513 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15430 \$153 \$11444 \$10370 \$11065 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15432 \$16 \$11399 \$16 \$153 \$11065 VNB sky130_fd_sc_hd__inv_1
X$15433 \$16 \$11399 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15434 \$16 \$10300 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15436 \$153 \$11376 \$11410 \$10386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15437 \$153 \$11478 \$11410 \$10300 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15438 \$16 \$10386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15439 \$153 \$11478 \$10417 \$11354 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15442 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$15443 \$16 \$10809 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15445 \$153 \$11642 \$11410 \$10809 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15446 \$16 \$10551 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15447 \$153 \$11540 \$11410 \$10551 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15448 \$16 \$12347 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15449 \$16 \$11013 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15450 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$15452 \$16 \$10578 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15453 \$16 \$10735 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15455 \$153 \$11445 \$11410 \$10735 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15456 \$153 \$11541 \$11410 \$10578 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15457 \$153 \$11445 \$10919 \$11354 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15458 \$16 \$11502 \$16 \$153 \$11354 VNB sky130_fd_sc_hd__inv_1
X$15459 \$16 \$11502 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15461 \$16 \$10386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15463 \$153 \$11379 \$11355 \$10386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15464 \$16 \$10551 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15466 \$153 \$11491 \$11355 \$10551 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15468 \$153 \$11491 \$10471 \$11215 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15470 \$16 \$10735 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15471 \$153 \$11356 \$11355 \$10735 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15472 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$15474 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$15475 \$153 \$11514 \$10714 \$11215 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15477 \$16 \$10300 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15478 \$16 \$10809 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15479 \$153 \$11446 \$11278 \$10300 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15480 \$16 \$10809 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15482 \$16 \$10551 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15483 \$153 \$11542 \$11278 \$10551 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15485 \$153 \$11309 \$10501 \$11215 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15487 \$16 \$10578 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15488 \$153 \$11411 \$11278 \$10578 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15489 \$153 \$11380 \$10919 \$10948 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15491 \$16 \$11496 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15492 \$153 \$11411 \$10370 \$10948 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15493 \$16 \$11496 \$16 \$153 \$10948 VNB sky130_fd_sc_hd__inv_1
X$15496 \$16 \$11496 \$11412 \$11543 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$15497 \$16 \$11412 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15498 \$16 \$10386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15499 \$153 \$11447 \$11279 \$10386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15500 \$16 \$10809 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15501 \$153 \$11544 \$11279 \$10809 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15502 \$16 \$11496 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15505 \$16 \$10611 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15506 \$16 \$11413 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15507 \$153 \$11545 \$11279 \$10611 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15509 \$153 \$11448 \$10417 \$11219 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15511 \$16 \$10578 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15512 \$153 \$11334 \$10501 \$11270 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15513 \$153 \$11447 \$10472 \$11219 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15514 \$153 \$11449 \$11311 \$10578 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15516 \$16 \$11546 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15517 \$16 \$10611 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15519 \$153 \$11547 \$11311 \$10611 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15520 \$153 \$11414 \$10501 \$11673 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15521 \$153 \$11479 \$11311 \$10735 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15522 \$153 \$11449 \$10370 \$11270 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15525 \$153 \$11450 \$11311 \$10551 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15526 \$153 \$11479 \$10919 \$11270 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15528 \$153 \$11311 \$11385 \$11492 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$15529 \$153 \$11450 \$10471 \$11270 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15530 \$16 \$7656 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15531 \$16 \$7656 \$16 \$153 \$11359 VNB sky130_fd_sc_hd__clkbuf_2
X$15533 \$16 \$11546 \$11412 \$11492 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$15535 \$16 \$10478 \$16 \$153 \$11358 VNB sky130_fd_sc_hd__clkbuf_2
X$15536 \$16 \$10478 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15537 \$153 \$11357 \$11359 \$11549 \$11358 \$16 \$16 VNB
+ sky130_fd_sc_hd__nor3b_4
X$15538 \$16 \$11357 \$11358 \$11359 \$153 \$11415 \$16 VNB
+ sky130_fd_sc_hd__and3b_4
X$15539 \$16 \$11415 \$16 \$153 \$11223 VNB sky130_fd_sc_hd__clkbuf_2
X$15540 \$16 \$11451 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15541 \$16 \$11383 \$16 \$153 \$10854 VNB sky130_fd_sc_hd__clkbuf_2
X$15542 \$16 \$11381 \$16 \$153 \$11374 VNB sky130_fd_sc_hd__clkbuf_2
X$15543 \$153 \$11503 \$10587 \$11016 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15545 \$16 \$11399 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15546 \$16 \$11382 \$16 \$153 \$11399 VNB sky130_fd_sc_hd__clkbuf_2
X$15547 \$153 \$11452 \$11451 \$11416 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$15548 \$153 \$11281 \$11578 \$11493 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$15549 \$16 \$11399 \$16 \$153 \$11226 VNB sky130_fd_sc_hd__inv_1
X$15550 \$16 \$11399 \$10838 \$11493 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$15551 \$153 \$11453 \$11281 \$10392 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15552 \$16 \$10564 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15554 \$153 \$11480 \$11452 \$10564 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15555 \$153 \$11453 \$10815 \$11226 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15556 \$153 \$11480 \$10642 \$11515 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15557 \$16 \$10564 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15558 \$16 \$10392 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15559 \$16 \$11016 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15560 \$16 \$11399 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15561 \$16 \$11016 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15562 \$16 \$11360 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15564 \$153 \$11454 \$11452 \$10346 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15565 \$16 \$11318 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15567 \$153 \$11481 \$11452 \$10617 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15568 \$16 \$10346 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15569 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$15570 \$16 \$10617 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15571 \$16 \$10393 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15573 \$153 \$11455 \$11281 \$10617 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15574 \$16 \$11502 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15577 \$16 \$11604 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15578 \$16 \$11502 \$11504 \$11494 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$15579 \$153 \$11316 \$11604 \$11494 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$15580 \$153 \$11455 \$10560 \$11226 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15581 \$16 \$10617 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15582 \$16 \$10617 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15583 \$153 \$11550 \$11316 \$10617 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15584 \$16 \$10446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15587 \$153 \$11227 \$11316 \$10446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15588 \$16 \$10393 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15589 \$153 \$11457 \$11316 \$10392 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15590 \$153 \$11456 \$11316 \$10326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15592 \$153 \$11550 \$10560 \$11384 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15593 \$153 \$11456 \$10466 \$11384 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15594 \$16 \$10446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15595 \$153 \$11552 \$11283 \$10446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15596 \$153 \$11457 \$10815 \$11384 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15597 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$15598 \$16 \$11622 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15600 \$16 \$11622 \$16 \$153 \$11495 VNB sky130_fd_sc_hd__inv_1
X$15601 \$16 \$10564 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15602 \$153 \$11482 \$11283 \$10564 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15604 \$16 \$10467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15605 \$153 \$11458 \$11283 \$10467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15607 \$153 \$11482 \$10642 \$11495 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15608 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$15610 \$16 \$10326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15612 \$153 \$11391 \$10560 \$11390 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15613 \$153 \$11458 \$10587 \$11495 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15614 \$153 \$11503 \$11346 \$10467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15615 \$16 \$11496 \$11229 \$11553 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$15616 \$16 \$10617 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15617 \$153 \$11554 \$11346 \$10617 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15618 \$16 \$11390 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15620 \$16 \$11496 \$16 \$153 \$11016 VNB sky130_fd_sc_hd__inv_1
X$15621 \$16 \$10564 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15623 \$153 \$11555 \$11346 \$10446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15624 \$153 \$11360 \$11346 \$10564 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15625 \$16 \$11459 \$11229 \$11497 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$15626 \$16 \$11459 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15627 \$16 \$11496 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15628 \$16 \$10393 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15629 \$16 \$11747 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15630 \$153 \$11460 \$11285 \$10393 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15632 \$153 \$11285 \$11747 \$11497 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$15634 \$153 \$10363 \$10466 \$10858 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15635 \$153 \$11517 \$11285 \$10564 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15636 \$16 \$10564 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15637 \$16 \$10467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15639 \$153 \$11392 \$11285 \$10467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15640 \$153 \$11021 \$10694 \$11516 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15641 \$16 \$10446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15642 \$153 \$11498 \$11385 \$11556 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$15643 \$16 \$10564 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15644 \$16 \$11946 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15645 \$153 \$11230 \$11946 \$11417 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$15647 \$16 \$11483 \$11229 \$11417 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$15648 \$153 \$11557 \$11498 \$10326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15649 \$153 \$13022 \$11498 \$10393 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15651 \$16 \$11546 \$16 \$153 \$12782 VNB sky130_fd_sc_hd__inv_1
X$15652 \$16 \$10564 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15653 \$16 \$11483 \$16 \$153 \$11461 VNB sky130_fd_sc_hd__inv_1
X$15654 \$153 \$10567 \$10694 \$10801 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15656 \$153 \$11462 \$11498 \$10564 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15657 \$153 \$11558 \$11498 \$10346 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15659 \$153 \$11463 \$11498 \$10392 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15660 \$16 \$10346 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15661 \$16 \$10392 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15662 \$16 \$11546 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15665 \$16 \$10467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15666 \$153 \$11559 \$11498 \$10467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15667 \$153 \$11464 \$11230 \$10392 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15669 \$153 \$10803 \$10587 \$10741 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15670 \$16 \$10392 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15671 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$15674 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$15675 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$15676 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$15677 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$15678 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$15679 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$15680 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$15681 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$15682 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$15683 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$15684 \$153 \$12511 \$12355 \$12294 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15687 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$15689 \$153 \$12638 \$12208 \$12512 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15690 \$16 \$12294 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15692 \$153 \$12561 \$12355 \$12236 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15694 \$153 \$12655 \$12656 \$12236 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15697 \$153 \$12561 \$12134 \$12386 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15698 \$16 \$12236 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15699 \$16 \$11078 \$16 \$153 \$12512 VNB sky130_fd_sc_hd__inv_1
X$15701 \$153 \$12656 \$11004 \$12584 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$15702 \$16 \$11078 \$12012 \$12584 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$15704 \$153 \$12438 \$12355 \$12095 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15705 \$16 \$12236 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15706 \$16 \$11004 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15708 \$16 \$12095 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15709 \$16 \$11078 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15710 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$15711 \$153 \$12585 \$12353 \$12512 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15712 \$153 \$12613 \$12134 \$12563 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15713 \$16 \$12095 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15714 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$15715 \$153 \$12613 \$12469 \$12236 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15716 \$153 \$12468 \$11810 \$12563 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15718 \$153 \$12562 \$12469 \$12095 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15720 \$153 \$12523 \$12229 \$12563 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15722 \$153 \$12562 \$12353 \$12563 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15723 \$16 \$12095 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15725 \$153 \$12614 \$12209 \$12563 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15726 \$153 \$12524 \$12057 \$12563 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15728 \$16 \$10939 \$16 \$153 \$12563 VNB sky130_fd_sc_hd__inv_1
X$15729 \$16 \$12152 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15732 \$153 \$12440 \$12586 \$12236 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15733 \$153 \$12586 \$10523 \$12525 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$15734 \$16 \$12564 \$16 \$153 \$12012 VNB sky130_fd_sc_hd__clkbuf_2
X$15735 \$153 \$12526 \$12353 \$12426 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15736 \$16 \$10523 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15739 \$153 \$12441 \$12586 \$12003 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15740 \$153 \$12639 \$12208 \$12426 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15742 \$153 \$12640 \$12412 \$12426 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15743 \$16 \$10453 \$16 \$153 \$12426 VNB sky130_fd_sc_hd__inv_1
X$15744 \$16 \$12003 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15746 \$16 \$12093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15747 \$16 \$10453 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15748 \$153 \$12587 \$12471 \$12093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15749 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$15751 \$153 \$12657 \$12471 \$12294 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15752 \$16 \$12294 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15753 \$153 \$12528 \$12353 \$12578 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15754 \$153 \$12587 \$12229 \$12578 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15756 \$16 \$12564 \$16 \$153 \$12015 VNB sky130_fd_sc_hd__clkbuf_2
X$15757 \$16 \$8361 \$16 \$153 \$12564 VNB sky130_fd_sc_hd__clkbuf_2
X$15759 \$153 \$12377 \$12471 \$12236 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15760 \$153 \$12658 \$12471 \$12230 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15761 \$16 \$11077 \$16 \$153 \$12578 VNB sky130_fd_sc_hd__inv_1
X$15762 \$153 \$12529 \$12057 \$12578 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15763 \$16 \$12236 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15765 \$153 \$12588 \$12444 \$12095 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15766 \$16 \$12230 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15768 \$16 \$11077 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15769 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$15770 \$153 \$12588 \$12353 \$12413 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15771 \$153 \$12589 \$12444 \$12158 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15772 \$153 \$12659 \$12444 \$12236 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15773 \$16 \$12158 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15775 \$16 \$12095 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15776 \$16 \$12236 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15777 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$15778 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$15779 \$16 \$10747 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15780 \$153 \$12590 \$12514 \$12158 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15781 \$153 \$12514 \$10624 \$12530 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$15782 \$16 \$10624 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15783 \$16 \$12158 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15785 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$15787 \$153 \$12495 \$12353 \$12579 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15789 \$153 \$12591 \$12514 \$12003 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15790 \$153 \$12590 \$12057 \$12579 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15791 \$16 \$12003 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15792 \$153 \$12496 \$12229 \$12579 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15793 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$15794 \$16 \$12158 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15795 \$153 \$12660 \$12391 \$12236 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15797 \$153 \$12592 \$12391 \$12158 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15798 \$16 \$12152 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15800 \$153 \$12531 \$12353 \$12392 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15801 \$153 \$12592 \$12057 \$12392 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15803 \$16 \$12236 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15804 \$153 \$12473 \$12229 \$12392 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15807 \$153 \$12532 \$12208 \$12392 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15808 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$15809 \$16 \$16 \$153 VNB sky130_fd_sc_hd__conb_1
X$15810 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$15811 \$16 \$11078 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15812 \$153 \$153 \$12208 \$12415 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15813 \$153 \$153 \$12229 \$12415 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15814 \$16 \$11004 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15815 \$153 \$12615 \$11004 \$12661 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$15816 \$16 \$10500 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15817 \$16 \$10888 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15819 \$153 \$153 \$12412 \$12415 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15820 \$16 \$10634 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15822 \$153 \$12616 \$12615 \$12296 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15824 \$153 \$12565 \$12357 \$12259 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15828 \$153 \$12616 \$12359 \$12641 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15829 \$153 \$12565 \$12307 \$12427 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15830 \$16 \$11078 \$16 \$153 \$12641 VNB sky130_fd_sc_hd__inv_1
X$15832 \$153 \$12515 \$12357 \$12083 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15833 \$16 \$12296 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15834 \$153 \$12642 \$12615 \$12160 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15836 \$16 \$12083 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15837 \$16 \$12160 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15838 \$153 \$12662 \$12533 \$12101 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15839 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$15840 \$153 \$12593 \$12533 \$12044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15841 \$153 \$12642 \$12028 \$12641 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15842 \$16 \$12044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15843 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$15846 \$153 \$12617 \$12533 \$12259 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15847 \$153 \$12594 \$12533 \$12295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15848 \$153 \$12535 \$12028 \$12154 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15849 \$153 \$12617 \$12307 \$12154 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15850 \$16 \$12295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15851 \$16 \$12259 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15853 \$16 \$12581 \$16 \$153 \$12159 VNB sky130_fd_sc_hd__clkbuf_2
X$15854 \$153 \$12710 \$10523 \$12536 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$15855 \$153 \$12618 \$12477 \$12241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15857 \$153 \$12499 \$12476 \$12498 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15858 \$153 \$12618 \$12363 \$12498 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15859 \$153 \$12447 \$12477 \$12160 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15861 \$153 \$12619 \$12068 \$12498 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15862 \$16 \$12241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15864 \$16 \$12160 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15865 \$153 \$12537 \$12174 \$12498 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15866 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$15867 \$153 \$12580 \$12710 \$12044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15868 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$15870 \$16 \$12044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15871 \$153 \$12580 \$12068 \$12729 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15873 \$153 \$12643 \$12476 \$12729 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15874 \$16 \$12581 \$16 \$153 \$12161 VNB sky130_fd_sc_hd__clkbuf_2
X$15875 \$16 \$11297 \$12161 \$12663 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$15876 \$153 \$12448 \$12500 \$12295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15877 \$153 \$12644 \$12359 \$12360 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15879 \$16 \$11297 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15880 \$16 \$12295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15881 \$16 \$7894 \$16 \$153 \$12581 VNB sky130_fd_sc_hd__clkbuf_2
X$15882 \$153 \$12645 \$12476 \$12758 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15884 \$153 \$12480 \$12500 \$12101 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15885 \$16 \$7894 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15887 \$153 \$12664 \$12500 \$12259 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15888 \$16 \$12101 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15891 \$153 \$12539 \$12174 \$12360 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15892 \$153 \$12620 \$12500 \$12044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15893 \$16 \$12259 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15895 \$153 \$12595 \$12508 \$12083 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15896 \$16 \$12044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15897 \$16 \$11077 \$16 \$153 \$12429 VNB sky130_fd_sc_hd__inv_1
X$15898 \$16 \$11077 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15901 \$153 \$12620 \$12068 \$12360 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15902 \$153 \$12595 \$12174 \$12429 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15903 \$16 \$12296 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15904 \$16 \$12083 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15905 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$15906 \$153 \$12566 \$12502 \$12259 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15907 \$153 \$12449 \$12502 \$12296 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15909 \$16 \$12259 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15910 \$16 \$12296 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15911 \$153 \$12733 \$12363 \$12429 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15912 \$153 \$12566 \$12307 \$12430 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15913 \$153 \$12450 \$12502 \$12101 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15915 \$16 \$12295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15917 \$16 \$11594 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15918 \$153 \$12541 \$12308 \$12296 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15921 \$16 \$12101 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15922 \$16 \$10974 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15923 \$16 \$12160 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15924 \$153 \$12665 \$12621 \$12160 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15925 \$16 \$12296 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15927 \$153 \$12567 \$12308 \$12160 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15928 \$153 \$12666 \$12621 \$12295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15929 \$16 \$12160 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15931 \$153 \$12567 \$12028 \$12378 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15933 \$16 \$12044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15934 \$16 \$12295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15935 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$15936 \$153 \$12667 \$12621 \$12044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15937 \$16 \$12241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15938 \$153 \$12596 \$12621 \$12241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15940 \$153 \$153 \$12363 \$12431 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15941 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$15943 \$153 \$12667 \$12068 \$12704 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15944 \$16 \$12115 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15945 \$153 \$12597 \$12400 \$12571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15947 \$16 \$12297 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15948 \$153 \$12622 \$12400 \$12297 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15950 \$153 \$12568 \$12400 \$12115 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15951 \$16 \$12297 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15952 \$153 \$12622 \$12582 \$12325 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15953 \$153 \$12568 \$12234 \$12325 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15955 \$16 \$10831 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15956 \$16 \$10831 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15957 \$16 \$12219 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15958 \$16 \$12233 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15959 \$153 \$12569 \$12400 \$12219 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15961 \$153 \$12516 \$12400 \$12233 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15962 \$153 \$12569 \$12110 \$12325 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15963 \$16 \$10831 \$12379 \$12668 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$15965 \$153 \$12623 \$12482 \$12297 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15966 \$16 \$11148 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15967 \$16 \$12406 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15970 \$16 \$12115 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15972 \$16 \$12326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15973 \$153 \$12481 \$12165 \$12517 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15974 \$153 \$12623 \$12582 \$12517 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15975 \$153 \$12598 \$12482 \$12326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15976 \$153 \$12646 \$12603 \$12517 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15978 \$153 \$12624 \$12482 \$12571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15979 \$153 \$12570 \$12482 \$12164 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15980 \$153 \$12598 \$12264 \$12517 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15981 \$153 \$12570 \$12217 \$12517 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15982 \$153 \$12624 \$12309 \$12517 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15984 \$16 \$10780 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15985 \$16 \$12219 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15986 \$153 \$12599 \$12518 \$12219 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15987 \$16 \$12600 \$16 \$153 \$12379 VNB sky130_fd_sc_hd__clkbuf_2
X$15988 \$153 \$12647 \$12582 \$12503 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15989 \$153 \$12599 \$12110 \$12503 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15990 \$16 \$8361 \$16 \$153 \$12600 VNB sky130_fd_sc_hd__clkbuf_2
X$15991 \$16 \$8361 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15993 \$153 \$12601 \$12518 \$12164 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$15995 \$153 \$12546 \$12264 \$12503 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15996 \$16 \$12164 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$15997 \$153 \$12601 \$12217 \$12503 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15998 \$153 \$12547 \$12234 \$12503 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$15999 \$153 \$12625 \$12165 \$12503 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16001 \$16 \$12164 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16003 \$153 \$12453 \$12452 \$12164 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16004 \$16 \$12600 \$16 \$153 \$12634 VNB sky130_fd_sc_hd__clkbuf_2
X$16005 \$16 \$11622 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16006 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$16007 \$16 \$12219 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16008 \$16 \$12571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16010 \$153 \$12454 \$12452 \$12571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16011 \$16 \$12612 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16012 \$153 \$12626 \$12165 \$12648 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16014 \$16 \$12233 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16015 \$153 \$12649 \$12110 \$12432 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16016 \$16 \$11622 \$16 \$153 \$12432 VNB sky130_fd_sc_hd__inv_1
X$16017 \$16 \$11622 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16018 \$16 \$12233 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16019 \$153 \$12602 \$12113 \$12233 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16020 \$16 \$12600 \$16 \$153 \$12166 VNB sky130_fd_sc_hd__clkbuf_2
X$16022 \$153 \$12669 \$12670 \$12164 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16024 \$153 \$12602 \$12603 \$12200 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16025 \$16 \$12164 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16026 \$153 \$12670 \$10615 \$12604 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$16027 \$16 \$10552 \$12166 \$12604 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$16029 \$16 \$12297 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16030 \$153 \$12572 \$12075 \$12297 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16031 \$16 \$12297 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16032 \$16 \$10615 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16033 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$16035 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$16036 \$153 \$12572 \$12582 \$11999 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16037 \$153 \$12504 \$12165 \$11999 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16038 \$153 \$12550 \$12309 \$11999 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16039 \$16 \$10552 \$16 \$153 \$12671 VNB sky130_fd_sc_hd__inv_1
X$16041 \$153 \$12627 \$12714 \$12164 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16042 \$16 \$12164 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16044 \$16 \$12326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16046 \$153 \$12456 \$12177 \$12326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16047 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$16049 \$153 \$12485 \$12309 \$12117 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16050 \$153 \$12551 \$12582 \$12117 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16051 \$153 \$12505 \$12165 \$12117 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16053 \$16 \$12297 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16055 \$153 \$12573 \$12204 \$12297 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16056 \$153 \$12672 \$12204 \$12298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16057 \$153 \$12573 \$12582 \$12333 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16059 \$16 \$12571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16060 \$153 \$12673 \$12605 \$12571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16062 \$16 \$12164 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16064 \$16 \$12115 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16065 \$153 \$12605 \$10960 \$12552 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$16066 \$153 \$12674 \$12605 \$12298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16067 \$153 \$12519 \$12204 \$12115 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16068 \$16 \$12233 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16069 \$16 \$12348 \$11776 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$16071 \$153 \$12628 \$12605 \$12233 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16072 \$153 \$12520 \$12204 \$12326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16073 \$153 \$12628 \$12603 \$12488 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16074 \$16 \$12433 \$12612 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$16075 \$16 \$10854 \$12459 \$12606 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$16077 \$153 \$12675 \$10780 \$12606 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$16079 \$16 \$12287 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16080 \$153 \$153 \$12182 \$12405 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16082 \$153 \$12629 \$12675 \$12287 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16083 \$153 \$153 \$11881 \$12405 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16084 \$153 \$153 \$12227 \$12405 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16086 \$153 \$12629 \$12339 \$12650 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16087 \$16 \$16 \$153 VNB sky130_fd_sc_hd__conb_1
X$16089 \$153 \$12607 \$12434 \$11983 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16091 \$153 \$12651 \$12119 \$12650 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16092 \$153 \$12607 \$11881 \$12423 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16093 \$16 \$11983 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16094 \$16 \$12351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16095 \$16 \$11113 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16097 \$16 \$10978 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16098 \$16 \$10831 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16100 \$16 \$10831 \$12459 \$12676 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$16101 \$153 \$12553 \$12371 \$12423 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16102 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$16103 \$16 \$12384 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16104 \$153 \$12608 \$12434 \$12384 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16105 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$16108 \$16 \$10831 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16109 \$153 \$12609 \$12434 \$12120 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16110 \$153 \$12608 \$12179 \$12423 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16111 \$153 \$12609 \$12182 \$12423 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16112 \$16 \$7894 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16113 \$16 \$12574 \$16 \$153 \$12459 VNB sky130_fd_sc_hd__clkbuf_2
X$16114 \$153 \$12630 \$12489 \$12287 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16115 \$16 \$7894 \$16 \$153 \$12574 VNB sky130_fd_sc_hd__clkbuf_2
X$16117 \$153 \$12383 \$12489 \$12351 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16118 \$16 \$12287 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16119 \$153 \$12761 \$12227 \$12337 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16121 \$153 \$12463 \$12489 \$12120 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16122 \$153 \$12630 \$12339 \$12337 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16125 \$16 \$12612 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16126 \$153 \$12583 \$12612 \$12677 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$16127 \$16 \$12120 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16128 \$153 \$12464 \$12583 \$12287 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16129 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$16130 \$16 \$12010 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16132 \$153 \$12652 \$12227 \$12435 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16133 \$16 \$12384 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16136 \$153 \$12466 \$12583 \$12010 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16137 \$153 \$12653 \$12119 \$12435 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16138 \$153 \$12124 \$12182 \$12147 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16139 \$16 \$10615 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16140 \$16 \$12574 \$16 \$153 \$12018 VNB sky130_fd_sc_hd__clkbuf_2
X$16141 \$153 \$12635 \$10615 \$12555 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$16142 \$16 \$12574 \$16 \$153 \$12678 VNB sky130_fd_sc_hd__clkbuf_2
X$16146 \$153 \$12679 \$12635 \$12351 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16147 \$16 \$12351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16148 \$16 \$12351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16149 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$16150 \$153 \$12556 \$12119 \$12302 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16151 \$16 \$10552 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16152 \$16 \$11983 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16153 \$16 \$10552 \$16 \$153 \$12680 VNB sky130_fd_sc_hd__inv_1
X$16154 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$16155 \$153 \$12681 \$12635 \$11983 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16158 \$16 \$12351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16159 \$153 \$12557 \$12179 \$12302 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16160 \$153 \$12631 \$12635 \$12384 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16161 \$16 \$12384 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16162 \$153 \$12610 \$12088 \$12351 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16164 \$153 \$12631 \$12179 \$12680 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16166 \$16 \$12120 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16167 \$153 \$12490 \$12339 \$12127 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16169 \$153 \$12682 \$12409 \$12120 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16170 \$153 \$12610 \$12119 \$12127 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16171 \$16 \$11983 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16172 \$16 \$12299 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16173 \$153 \$12632 \$12409 \$12299 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16176 \$153 \$12611 \$11881 \$12521 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16178 \$153 \$12575 \$12409 \$12010 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16180 \$153 \$12632 \$12371 \$12521 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16181 \$16 \$11280 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16182 \$153 \$12575 \$11942 \$12521 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16183 \$16 \$11385 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16185 \$16 \$11983 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16186 \$153 \$12683 \$12636 \$11983 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16188 \$16 \$11546 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16189 \$16 \$12287 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16190 \$153 \$12576 \$12373 \$12287 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16191 \$153 \$12637 \$12636 \$12287 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16193 \$153 \$12576 \$12339 \$12411 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16194 \$16 \$12351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16195 \$16 \$12299 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16196 \$153 \$11323 \$10560 \$11322 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16197 \$153 \$12684 \$12636 \$12299 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16198 \$153 \$12577 \$12373 \$12351 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16199 \$16 \$12384 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16201 \$153 \$12633 \$12636 \$12384 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16202 \$153 \$12577 \$12119 \$12411 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16203 \$153 \$11792 \$10466 \$11926 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16204 \$153 \$12684 \$12371 \$12654 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16205 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$16206 \$153 \$12637 \$12339 \$12654 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16208 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$16209 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$16210 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$16211 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$16212 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$16213 \$153 \$3284 \$2006 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$16214 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$16215 \$153 \$3390 \$3389 \$3208 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16216 \$153 \$3391 \$3606 \$3208 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16217 \$153 \$3285 \$3207 \$2006 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16219 \$153 \$3445 \$3478 \$3208 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16221 \$153 \$3066 \$3207 \$1942 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16222 \$153 \$3550 \$3394 \$3420 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16223 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$16225 \$153 \$3067 \$3207 \$2024 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16226 \$16 \$1942 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16228 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$16230 \$153 \$3214 \$3207 \$2180 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16231 \$153 \$3421 \$3422 \$3420 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16232 \$16 \$2180 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16233 \$16 \$3571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16234 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$16235 \$16 \$2024 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16236 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$16239 \$153 \$3287 \$3170 \$1687 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16240 \$153 \$3392 \$3170 \$2024 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16241 \$153 \$3330 \$3394 \$3331 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16242 \$153 \$3423 \$3540 \$3331 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16243 \$16 \$1687 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16244 \$153 \$3424 \$3307 \$3331 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16247 \$153 \$3215 \$3170 \$2180 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16249 \$153 \$3446 \$3497 \$3385 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16250 \$153 \$3332 \$3170 \$1795 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16251 \$16 \$3385 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16252 \$16 \$3473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16255 \$153 \$3425 \$3422 \$3426 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16256 \$16 \$2180 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16257 \$16 \$1795 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16258 \$16 \$1404 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16259 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$16261 \$153 \$3300 \$3148 \$1942 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16262 \$153 \$3393 \$3407 \$3571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16264 \$153 \$3332 \$1815 \$3056 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16265 \$153 \$3393 \$3422 \$3578 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16266 \$153 \$3299 \$1547 \$3056 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16267 \$153 \$3427 \$3394 \$3578 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16268 \$153 \$3197 \$3148 \$1795 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16269 \$16 \$3571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16270 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$16272 \$153 \$3428 \$3490 \$3578 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16273 \$153 \$3301 \$2210 \$3149 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16274 \$16 \$1795 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16275 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$16276 \$153 \$3300 \$2064 \$3149 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16278 \$153 \$3447 \$3408 \$3571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16279 \$16 \$1594 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16280 \$16 \$1942 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16282 \$153 \$3345 \$3093 \$2024 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16283 \$16 \$3571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16284 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$16285 \$153 \$3429 \$3394 \$3476 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16286 \$16 \$2024 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16287 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$16288 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$16289 \$153 \$3333 \$1687 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$16292 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$16293 \$153 \$3430 \$3540 \$3409 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16294 \$153 \$3345 \$2210 \$3015 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16295 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$16296 \$153 \$3431 \$3394 \$3409 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16297 \$16 \$3333 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16298 \$16 \$1551 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16300 \$16 \$3474 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16302 \$153 \$3304 \$3017 \$2024 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16304 \$153 \$3396 \$3410 \$3615 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16305 \$16 \$2024 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16307 \$153 \$3346 \$3394 \$3334 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16308 \$153 \$3395 \$3490 \$3334 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16311 \$153 \$3396 \$3307 \$3334 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16312 \$153 \$3335 \$1942 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$16313 \$16 \$3615 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16314 \$16 \$1508 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16315 \$16 \$1332 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16316 \$16 \$2743 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16317 \$153 \$1406 \$3571 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$16318 \$16 \$3335 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16320 \$16 \$2743 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16321 \$16 \$2064 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16324 \$16 \$1406 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16325 \$153 \$3244 \$1658 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$16327 \$16 \$1625 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16328 \$153 \$3448 \$1482 \$2064 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16329 \$16 \$3244 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16331 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16333 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16334 \$153 \$3449 \$1482 \$2252 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16335 \$153 \$3365 \$1482 \$1792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16336 \$153 \$3397 \$1482 \$2210 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16337 \$153 \$153 \$1547 \$3151 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16340 \$153 \$3305 \$1482 \$3490 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16341 \$153 \$3450 \$1482 \$1547 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16342 \$153 \$3366 \$1482 \$3422 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16343 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16344 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16345 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16346 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16348 \$153 \$3239 \$1482 \$3394 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16349 \$16 \$3540 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16350 \$16 \$3422 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16351 \$153 \$3367 \$3005 \$1965 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16352 \$16 \$3394 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16353 \$16 \$2210 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16355 \$153 \$3451 \$3412 \$3573 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16356 \$16 \$1965 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16357 \$16 \$1496 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16359 \$16 \$1508 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16361 \$16 \$3573 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16362 \$153 \$3368 \$3005 \$2042 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16363 \$153 \$3367 \$1806 \$3269 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16364 \$153 \$3368 \$1924 \$3269 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16365 \$16 \$2042 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16366 \$16 \$3555 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16368 \$153 \$3290 \$3005 \$2043 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16371 \$153 \$3347 \$3412 \$3492 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16372 \$153 \$3347 \$3354 \$3336 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16373 \$153 \$3432 \$3435 \$3336 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16374 \$16 \$2043 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16376 \$16 \$3492 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16377 \$16 \$1208 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16378 \$153 \$3398 \$3713 \$3573 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16380 \$153 \$3043 \$3144 \$2042 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16381 \$153 \$3398 \$3079 \$3583 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16382 \$16 \$3573 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16383 \$16 \$2042 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16385 \$153 \$3075 \$3144 \$1965 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16386 \$16 \$3386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16389 \$153 \$3260 \$2026 \$2879 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16391 \$153 \$3348 \$3354 \$3337 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16392 \$16 \$1965 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16394 \$153 \$3349 \$3502 \$3386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16395 \$153 \$3338 \$3079 \$3337 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16397 \$153 \$3349 \$3435 \$3337 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16399 \$153 \$3399 \$3413 \$3386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16400 \$16 \$3386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16401 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$16402 \$153 \$3350 \$3354 \$3339 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16403 \$153 \$3399 \$3435 \$3339 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16404 \$16 \$5596 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16405 \$16 \$3386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16406 \$16 \$1692 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16408 \$16 \$1750 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16409 \$153 \$3370 \$3309 \$1692 \$3414 \$5596 \$2075 \$3277 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$16410 \$153 \$3370 \$3369 \$1750 \$3257 \$3351 \$1664 \$3277 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$16411 \$153 \$3370 \$3416 \$1735 \$3479 \$3415 \$2407 \$3277 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$16412 \$16 \$3479 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16413 \$16 \$1735 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16416 \$16 \$3492 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16418 \$16 \$3307 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16419 \$153 \$3370 \$3371 \$1802 \$3557 \$3352 \$1925 \$3277 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$16420 \$16 \$3310 \$16 \$153 \$3370 VNB sky130_fd_sc_hd__clkbuf_2
X$16422 \$16 \$3270 \$3400 \$3371 \$235 \$16 \$153 VNB sky130_fd_sc_hd__mux2_1
X$16423 \$16 \$3241 \$16 \$153 \$3277 VNB sky130_fd_sc_hd__clkbuf_2
X$16425 \$153 \$3370 \$3452 \$1635 \$3481 \$3417 \$1597 \$3277 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$16426 \$153 \$3370 \$3372 \$1573 \$3239 \$3343 \$1294 \$3277 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$16427 \$16 \$3418 \$16 \$153 \$3270 VNB sky130_fd_sc_hd__clkbuf_2
X$16428 \$16 \$3239 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16429 \$16 \$1573 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16430 \$16 \$3418 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16432 \$16 \$1635 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16434 \$16 \$2364 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16435 \$153 \$3433 \$3079 \$3340 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16437 \$153 \$3220 \$3024 \$2043 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16438 \$16 \$3343 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16439 \$16 \$3417 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16440 \$16 \$3400 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16441 \$153 \$3434 \$3435 \$3340 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16442 \$153 \$3353 \$3354 \$3340 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16443 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$16444 \$16 \$2043 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16446 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$16447 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$16448 \$153 \$3291 \$3077 \$2042 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16449 \$153 \$3482 \$3504 \$3436 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16450 \$153 \$3453 \$3574 \$3386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16451 \$16 \$2042 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16453 \$16 \$3344 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16454 \$16 \$1965 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16456 \$153 \$3355 \$3077 \$1965 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16457 \$153 \$3437 \$3354 \$3436 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16458 \$153 \$3401 \$3079 \$3436 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16459 \$16 \$3310 \$3344 \$3241 \$153 \$1354 \$16 VNB sky130_fd_sc_hd__and3b_4
X$16460 \$153 \$153 \$1924 \$3292 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16461 \$16 \$1354 \$16 \$153 \$3292 VNB sky130_fd_sc_hd__clkbuf_2
X$16463 \$153 \$153 \$2026 \$3292 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16464 \$153 \$3439 \$1923 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$16465 \$153 \$153 \$1703 \$3292 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16466 \$16 \$3587 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16467 \$153 \$3587 \$1965 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$16468 \$16 \$3373 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16469 \$16 \$3439 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16470 \$16 \$3284 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16472 \$153 \$3355 \$1806 \$2908 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16474 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16475 \$153 \$3402 \$1482 \$2184 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16476 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16478 \$153 \$3284 \$2104 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$16480 \$153 \$3688 \$1482 \$1806 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16481 \$153 \$3244 \$1879 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$16482 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16486 \$153 \$3387 \$1482 \$3101 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16487 \$153 \$3333 \$1878 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$16488 \$16 \$3241 \$3344 \$3310 \$153 \$1378 \$16 VNB sky130_fd_sc_hd__and3b_4
X$16490 \$153 \$3127 \$3374 \$1705 \$3356 \$3357 \$1665 \$3139 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$16491 \$16 \$3310 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16494 \$16 \$3272 \$3454 \$3374 \$298 \$16 \$153 VNB sky130_fd_sc_hd__mux2_1
X$16495 \$153 \$3403 \$3281 \$1879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16496 \$16 \$3310 \$16 \$153 \$3127 VNB sky130_fd_sc_hd__clkbuf_2
X$16498 \$153 \$3313 \$1613 \$3341 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16499 \$153 \$3403 \$1558 \$3341 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16501 \$153 \$3127 \$3081 \$1706 \$3387 \$3358 \$3109 \$3139 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$16502 \$153 \$3455 \$3281 \$2098 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16504 \$153 \$3281 \$1628 \$3245 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$16505 \$16 \$3418 \$16 \$153 \$3272 VNB sky130_fd_sc_hd__clkbuf_2
X$16508 \$16 \$1566 \$16 \$153 \$3341 VNB sky130_fd_sc_hd__inv_1
X$16510 \$153 \$3294 \$3211 \$2104 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16511 \$16 \$1969 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16512 \$16 \$2098 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16513 \$153 \$3375 \$3211 \$2098 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16514 \$153 \$3455 \$1993 \$3341 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16516 \$16 \$3109 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16517 \$16 \$2935 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16519 \$153 \$3275 \$1558 \$3246 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16520 \$16 \$1756 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16521 \$153 \$3359 \$3282 \$1756 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16522 \$153 \$3359 \$1712 \$3246 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16523 \$16 \$2105 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16524 \$153 \$3314 \$2092 \$3246 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16525 \$16 \$1566 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16526 \$16 \$1585 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16529 \$153 \$3484 \$1868 \$3246 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16530 \$16 \$1708 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16531 \$16 \$1518 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16532 \$153 \$3315 \$1993 \$3246 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16533 \$16 \$3146 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16534 \$16 \$3103 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16535 \$16 \$3454 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16536 \$153 \$3247 \$1613 \$3246 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16537 \$16 \$2104 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16538 \$153 \$3404 \$3140 \$2104 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16539 \$16 \$3272 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16540 \$16 \$1879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16542 \$153 \$3224 \$3140 \$1879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16544 \$153 \$3404 \$2092 \$3162 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16546 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$16547 \$16 \$1756 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16548 \$153 \$3179 \$1613 \$3317 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16550 \$16 \$2104 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16551 \$153 \$3316 \$3225 \$2104 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16553 \$153 \$3405 \$3225 \$1756 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16555 \$153 \$3316 \$2092 \$3317 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16556 \$16 \$1879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16557 \$153 \$3457 \$3225 \$1879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16558 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$16561 \$16 \$1758 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16563 \$16 \$1969 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16564 \$153 \$3360 \$3283 \$1969 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16566 \$153 \$3361 \$3283 \$1756 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16567 \$16 \$2935 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16568 \$153 \$3361 \$1712 \$3131 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16569 \$16 \$1756 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16570 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$16572 \$153 \$3438 \$1715 \$3131 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16573 \$16 \$1599 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16574 \$153 \$3319 \$1993 \$3131 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16575 \$153 \$3457 \$1558 \$3317 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16576 \$153 \$3360 \$1613 \$3131 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16577 \$153 \$3458 \$3322 \$2104 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16578 \$16 \$2104 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16579 \$16 \$2016 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16581 \$16 \$1475 \$2935 \$3321 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$16582 \$153 \$3320 \$1993 \$3296 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16584 \$153 \$3297 \$3322 \$2016 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16585 \$153 \$3295 \$3322 \$1878 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16587 \$16 \$4223 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16588 \$16 \$3483 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16590 \$16 \$3456 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16591 \$16 \$2105 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16593 \$16 \$4414 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16594 \$153 \$3388 \$3322 \$2105 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16595 \$16 \$1879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16596 \$16 \$1756 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16597 \$153 \$3376 \$3322 \$1756 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16598 \$153 \$3228 \$3322 \$1879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16599 \$16 \$3402 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16601 \$153 \$3388 \$2438 \$3296 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16602 \$16 \$4408 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16605 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16606 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16607 \$153 \$3459 \$1482 \$2056 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16608 \$153 \$3377 \$1482 \$2267 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16609 \$16 \$2267 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16611 \$16 \$2056 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16612 \$16 \$393 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16614 \$16 \$1936 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16615 \$16 \$1475 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16616 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16617 \$16 \$1378 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16618 \$153 \$3199 \$2031 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$16619 \$153 \$3439 \$2085 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$16620 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16622 \$16 \$3199 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16623 \$16 \$3439 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16624 \$16 \$2085 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16625 \$16 \$2269 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16626 \$153 \$3378 \$3185 \$2085 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16628 \$153 \$3460 \$3185 \$2093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16629 \$153 \$3362 \$3185 \$2192 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16630 \$16 \$2093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16631 \$16 \$3461 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16632 \$16 \$3461 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16634 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$16636 \$153 \$3364 \$3185 \$1960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16637 \$153 \$3362 \$2269 \$3186 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16638 \$16 \$2192 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16639 \$153 \$3363 \$2000 \$3186 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16640 \$16 \$1960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16641 \$16 \$2093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16642 \$153 \$3406 \$3212 \$2093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16644 \$153 \$3364 \$2086 \$3186 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16645 \$16 \$1973 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16647 \$16 \$2085 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16648 \$153 \$3406 \$2265 \$3167 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16649 \$153 \$3379 \$3212 \$2085 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16650 \$16 \$2192 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16651 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$16654 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$16655 \$16 \$1860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16656 \$153 \$3440 \$2086 \$3167 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16657 \$16 \$1628 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16659 \$153 \$3323 \$1936 \$3342 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16660 \$153 \$3463 \$3250 \$1860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16661 \$153 \$2873 \$2000 \$2780 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16663 \$16 \$1566 \$16 \$153 \$3342 VNB sky130_fd_sc_hd__inv_1
X$16664 \$16 \$1566 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16665 \$16 \$1973 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16666 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$16667 \$153 \$3325 \$3250 \$1973 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16668 \$16 \$2192 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16669 \$153 \$3464 \$3250 \$2192 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16670 \$153 \$3133 \$2271 \$2780 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16671 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$16673 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$16674 \$153 \$2987 \$1936 \$2780 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16675 \$16 \$1860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16676 \$153 \$3465 \$3147 \$1860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16678 \$153 \$3380 \$3147 \$2031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16679 \$153 \$3466 \$3147 \$2085 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16681 \$153 \$3325 \$2056 \$3342 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16684 \$16 \$2093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16685 \$16 \$2192 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16686 \$153 \$3467 \$3251 \$2192 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16687 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$16688 \$16 \$2085 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16689 \$153 \$3143 \$3251 \$2085 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16691 \$153 \$3468 \$3251 \$2031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16692 \$16 \$1960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16693 \$16 \$2031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16695 \$16 \$2031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16696 \$153 \$3381 \$3252 \$2031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16697 \$153 \$3441 \$2086 \$2931 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16699 \$153 \$3381 \$1936 \$3169 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16701 \$153 \$3327 \$3252 \$2085 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16702 \$153 \$3469 \$3252 \$2192 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16703 \$153 \$3327 \$2271 \$3169 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16704 \$16 \$2192 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16705 \$16 \$1475 \$2984 \$3231 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$16706 \$16 \$1627 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16709 \$16 \$2984 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16710 \$16 \$2085 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16711 \$16 \$1758 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16712 \$153 \$3233 \$3253 \$2085 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16714 \$16 \$2085 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16715 \$153 \$3470 \$3254 \$2085 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16716 \$16 \$1758 \$16 \$153 \$3206 VNB sky130_fd_sc_hd__inv_1
X$16717 \$16 \$1475 \$16 \$153 \$3328 VNB sky130_fd_sc_hd__inv_1
X$16718 \$153 \$3442 \$2265 \$3206 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16719 \$16 \$2191 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16721 \$16 \$1758 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16722 \$16 \$1475 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16724 \$16 \$1973 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16725 \$153 \$3329 \$2267 \$3328 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16726 \$153 \$3382 \$3254 \$1973 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16727 \$153 \$3443 \$2265 \$3328 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16728 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$16729 \$16 \$2192 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16731 \$16 \$2031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16733 \$16 \$1960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16736 \$153 \$3383 \$3254 \$1960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16737 \$153 \$3471 \$3254 \$2031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16738 \$16 \$2031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16739 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$16740 \$153 \$3035 \$1936 \$2642 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16742 \$153 \$3444 \$2269 \$3206 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16744 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$16745 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$16746 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$16747 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$16748 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$16749 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$16750 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$16751 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$16752 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$16753 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$16756 \$153 \$12040 \$12019 \$12230 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16757 \$153 \$12040 \$12412 \$12020 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16759 \$153 \$12090 \$12019 \$12158 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16760 \$16 \$12230 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16761 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$16762 \$153 \$11959 \$10088 \$11717 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16764 \$153 \$12091 \$12019 \$12095 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16765 \$16 \$12158 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16767 \$16 \$11757 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16768 \$16 \$11987 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16770 \$153 \$11733 \$11987 \$11885 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$16771 \$16 \$12095 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16772 \$16 \$10348 \$12012 \$12130 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$16773 \$153 \$12021 \$12019 \$12003 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16774 \$16 \$10348 \$16 \$153 \$12020 VNB sky130_fd_sc_hd__inv_1
X$16775 \$16 \$10226 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16776 \$153 \$11988 \$11751 \$10226 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16779 \$153 \$11960 \$10088 \$11718 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16780 \$153 \$11988 \$10161 \$11718 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16782 \$16 \$11898 \$11347 \$12056 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$16783 \$16 \$10226 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16784 \$153 \$12092 \$12041 \$12095 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16786 \$153 \$11832 \$10276 \$11718 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16788 \$153 \$12021 \$11810 \$12020 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16789 \$153 \$12063 \$12041 \$12093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16790 \$153 \$12041 \$10522 \$12022 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$16791 \$16 \$10200 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16793 \$16 \$10539 \$16 \$153 \$12252 VNB sky130_fd_sc_hd__inv_1
X$16794 \$16 \$10539 \$12012 \$12022 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$16795 \$16 \$12158 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16797 \$153 \$11989 \$10890 \$12023 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$16798 \$153 \$12064 \$11810 \$12094 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16799 \$153 \$12064 \$11989 \$12003 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16800 \$153 \$11632 \$12013 \$11961 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$16801 \$153 \$12065 \$11989 \$12158 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16803 \$153 \$11990 \$11632 \$10200 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16804 \$153 \$12065 \$12057 \$12094 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16805 \$153 \$11990 \$10088 \$11560 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16806 \$16 \$10744 \$16 \$153 \$12094 VNB sky130_fd_sc_hd__inv_1
X$16807 \$16 \$10200 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16809 \$16 \$12095 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16810 \$153 \$11991 \$12014 \$12003 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16812 \$153 \$12066 \$12014 \$12095 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16813 \$153 \$11991 \$11810 \$12004 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16814 \$153 \$12066 \$12353 \$12004 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16815 \$16 \$12003 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16816 \$16 \$10367 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16818 \$153 \$12014 \$10722 \$12042 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$16820 \$153 \$11933 \$10330 \$11652 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16821 \$16 \$10555 \$12015 \$12042 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$16822 \$16 \$12093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16823 \$153 \$11892 \$10161 \$11652 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16824 \$153 \$12096 \$10706 \$12133 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$16825 \$153 \$12342 \$12134 \$12005 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16827 \$16 \$10722 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16828 \$16 \$10706 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16829 \$153 \$11992 \$11735 \$10200 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16831 \$16 \$12095 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16832 \$153 \$12024 \$12096 \$12158 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16833 \$16 \$10226 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16834 \$16 \$10200 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16835 \$16 \$12158 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16836 \$153 \$12097 \$12096 \$12003 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16837 \$16 \$11814 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16839 \$153 \$12024 \$12057 \$12005 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16840 \$16 \$11795 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16841 \$16 \$12003 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16843 \$153 \$12172 \$10667 \$12043 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$16844 \$16 \$10621 \$12015 \$12043 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$16845 \$16 \$10621 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16846 \$16 \$11995 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16847 \$153 \$12210 \$12229 \$12006 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16848 \$16 \$10667 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16850 \$153 \$12098 \$12353 \$12006 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16852 \$16 \$11814 \$11238 \$12025 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$16853 \$153 \$11801 \$12190 \$12025 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$16854 \$153 \$12099 \$12134 \$12006 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16856 \$153 \$8301 \$12158 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$16857 \$16 \$12190 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16858 \$16 \$11994 \$10682 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$16861 \$16 \$11994 \$11993 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$16862 \$153 \$11963 \$10088 \$11655 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16863 \$16 \$8301 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16864 \$16 \$11994 \$10722 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$16865 \$16 \$12016 \$11949 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$16866 \$16 \$11994 \$11364 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$16867 \$16 \$12016 \$12013 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$16868 \$16 \$12016 \$11190 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$16869 \$16 \$11943 \$16 \$153 \$12016 VNB sky130_fd_sc_hd__clkbuf_2
X$16870 \$16 \$12016 \$11432 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$16871 \$16 \$12016 \$11987 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$16872 \$16 \$12016 \$11567 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$16873 \$16 \$11994 \$11194 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$16875 \$16 \$11944 \$10634 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$16877 \$16 \$11805 \$11995 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$16878 \$16 \$11944 \$10603 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$16879 \$16 \$11805 \$11637 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$16880 \$16 \$11944 \$11004 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$16881 \$16 \$11805 \$11431 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$16882 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16884 \$153 \$10357 \$8340 \$11810 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16885 \$153 \$10165 \$8340 \$12209 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16887 \$16 \$10348 \$12159 \$12082 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$16888 \$16 \$11805 \$10959 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$16890 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16891 \$16 \$12209 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16892 \$153 \$10261 \$8340 \$12412 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16893 \$16 \$11810 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16894 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16895 \$153 \$10166 \$8340 \$12353 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16896 \$16 \$12412 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16898 \$16 \$12229 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16899 \$16 \$12353 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16900 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16902 \$153 \$12100 \$12191 \$12044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16903 \$153 \$10215 \$8340 \$12229 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16905 \$16 \$12044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16906 \$153 \$12102 \$12191 \$12083 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16907 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$16909 \$16 \$10522 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16910 \$16 \$10606 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16912 \$153 \$11964 \$10516 \$11818 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16913 \$153 \$12103 \$12191 \$12101 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16914 \$153 \$11996 \$10522 \$12026 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$16915 \$16 \$11757 \$11275 \$11965 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$16916 \$153 \$11997 \$11657 \$10605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16917 \$16 \$12101 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16919 \$153 \$12067 \$11996 \$12044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16920 \$153 \$11997 \$10686 \$11838 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16921 \$153 \$12067 \$12068 \$12238 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16922 \$16 \$10605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16924 \$16 \$11794 \$11275 \$11966 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$16925 \$16 \$12044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16926 \$153 \$12070 \$10890 \$12069 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$16929 \$153 \$11967 \$12013 \$11900 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$16930 \$16 \$10744 \$12159 \$12069 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$16931 \$153 \$11874 \$11658 \$10526 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16933 \$153 \$12105 \$12028 \$12104 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16935 \$16 \$10744 \$16 \$153 \$12104 VNB sky130_fd_sc_hd__inv_1
X$16936 \$16 \$10526 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16938 \$153 \$12106 \$12070 \$12083 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16939 \$16 \$10744 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16941 \$153 \$11950 \$11658 \$10605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16942 \$153 \$12084 \$10722 \$12138 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$16943 \$16 \$10605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16944 \$16 \$11721 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16947 \$16 \$10605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16948 \$153 \$12045 \$11967 \$10605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16949 \$153 \$12107 \$12084 \$12160 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16950 \$153 \$11877 \$11967 \$10606 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16951 \$16 \$10555 \$16 \$153 \$12071 VNB sky130_fd_sc_hd__inv_1
X$16952 \$16 \$12083 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16955 \$16 \$12160 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16956 \$16 \$10621 \$12161 \$12058 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$16957 \$16 \$10606 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16958 \$153 \$12027 \$12085 \$12101 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16959 \$153 \$12085 \$10667 \$12058 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$16961 \$16 \$12101 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16962 \$153 \$12059 \$12085 \$12160 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16963 \$16 \$10667 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16965 \$153 \$12027 \$12476 \$12007 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16966 \$16 \$10605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16967 \$16 \$12160 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16968 \$153 \$12108 \$12085 \$12083 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16970 \$153 \$12059 \$12028 \$12007 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16972 \$16 \$10413 \$12161 \$12046 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$16975 \$16 \$12083 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16976 \$153 \$12029 \$12068 \$12007 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16978 \$153 \$12086 \$10706 \$12046 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$16979 \$153 \$11902 \$10516 \$11488 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16980 \$153 \$11878 \$12086 \$12083 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16981 \$153 \$12030 \$12476 \$11869 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$16983 \$16 \$10470 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16985 \$16 \$10606 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16986 \$153 \$11952 \$11739 \$10606 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16987 \$16 \$10413 \$16 \$153 \$11869 VNB sky130_fd_sc_hd__inv_1
X$16989 \$153 \$12109 \$12086 \$12044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$16991 \$153 \$11806 \$12190 \$11969 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$16992 \$16 \$12044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$16996 \$153 \$8416 \$12160 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$16997 \$153 \$8734 \$12101 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$16998 \$153 \$11841 \$10401 \$11906 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17000 \$153 \$10311 \$12083 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$17001 \$153 \$10361 \$12044 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$17002 \$153 \$8821 \$8340 \$12028 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17003 \$16 \$10311 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17004 \$16 \$10361 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17005 \$16 \$9747 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17008 \$16 \$9138 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17009 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17010 \$153 \$9138 \$12164 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$17011 \$16 \$12028 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17012 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17013 \$153 \$8524 \$8340 \$12174 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17014 \$153 \$12072 \$10686 \$11906 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17016 \$16 \$12174 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17017 \$16 \$12155 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17018 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17019 \$16 \$8301 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17020 \$153 \$10180 \$8340 \$12234 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17021 \$153 \$8301 \$12219 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$17022 \$16 \$12582 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17023 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17024 \$153 \$11971 \$10370 \$11724 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17026 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17027 \$153 \$10322 \$8340 \$12110 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17028 \$153 \$10122 \$8340 \$12165 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17029 \$153 \$12111 \$11641 \$10300 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17030 \$16 \$11824 \$16 \$153 \$11724 VNB sky130_fd_sc_hd__inv_1
X$17031 \$16 \$10578 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17033 \$153 \$12047 \$11641 \$10578 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17035 \$16 \$12307 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17036 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17037 \$153 \$12047 \$10370 \$11665 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17038 \$153 \$12031 \$11641 \$10386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17039 \$16 \$10386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17041 \$16 \$12219 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17042 \$16 \$11930 \$16 \$153 \$11665 VNB sky130_fd_sc_hd__inv_1
X$17044 \$153 \$12111 \$10417 \$11665 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17045 \$153 \$12031 \$10472 \$11665 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17046 \$16 \$12115 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17047 \$16 \$11824 \$11378 \$12073 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$17049 \$153 \$11641 \$11842 \$12008 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$17050 \$153 \$11741 \$12162 \$12073 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$17052 \$153 \$11666 \$12009 \$11974 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$17053 \$153 \$11973 \$10501 \$11513 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17055 \$153 \$12033 \$11742 \$10300 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17057 \$16 \$12032 \$11378 \$12048 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$17058 \$153 \$11975 \$10472 \$11669 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17060 \$153 \$12033 \$10417 \$11669 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17061 \$153 \$12060 \$11742 \$10578 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17062 \$153 \$12060 \$10370 \$11669 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17064 \$153 \$12034 \$11880 \$10386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17065 \$16 \$12032 \$16 \$153 \$11669 VNB sky130_fd_sc_hd__inv_1
X$17066 \$16 \$10809 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17067 \$16 \$10386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17068 \$16 \$12032 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17071 \$16 \$10578 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17072 \$153 \$12034 \$10472 \$11725 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17073 \$16 \$11945 \$11378 \$12112 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$17074 \$153 \$12074 \$11880 \$10300 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17076 \$153 \$11998 \$11880 \$10578 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17077 \$16 \$10300 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17079 \$153 \$11998 \$10370 \$11725 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17080 \$153 \$12074 \$10417 \$11725 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17082 \$16 \$10736 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17083 \$153 \$12113 \$10981 \$12140 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$17085 \$16 \$10661 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17086 \$16 \$10981 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17087 \$16 \$10736 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17088 \$153 \$11911 \$10417 \$11954 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17089 \$153 \$11976 \$10472 \$11954 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17091 \$153 \$11807 \$11776 \$11912 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$17092 \$153 \$12114 \$12110 \$12200 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17093 \$153 \$11845 \$10501 \$11954 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17095 \$153 \$11775 \$10833 \$11954 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17096 \$16 \$10386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17097 \$16 \$12115 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17098 \$153 \$12049 \$11645 \$10386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17099 \$16 \$10661 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17101 \$16 \$12219 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17102 \$153 \$12075 \$12050 \$12116 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$17103 \$16 \$10649 \$16 \$153 \$11999 VNB sky130_fd_sc_hd__inv_1
X$17104 \$153 \$11977 \$10417 \$11727 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17105 \$153 \$8073 \$8340 \$12371 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17106 \$16 \$12050 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17109 \$16 \$10649 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17111 \$16 \$11798 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17112 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17113 \$153 \$11978 \$10370 \$11727 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17114 \$16 \$12371 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17116 \$153 \$12221 \$12110 \$12117 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17118 \$16 \$10578 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17119 \$153 \$12051 \$11808 \$10578 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17120 \$16 \$11798 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17121 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$17122 \$16 \$10853 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17125 \$16 \$11921 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17126 \$16 \$12219 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17127 \$153 \$11863 \$11808 \$10386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17129 \$153 \$12051 \$10370 \$11825 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17130 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$17131 \$16 \$10300 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17132 \$153 \$12076 \$11808 \$10300 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17133 \$16 \$10386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17134 \$16 \$11946 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17136 \$16 \$10809 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17138 \$153 \$11955 \$11808 \$10809 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17139 \$153 \$12118 \$10860 \$12205 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$17140 \$153 \$12076 \$10417 \$11825 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17141 \$16 \$10529 \$16 \$153 \$12246 VNB sky130_fd_sc_hd__inv_1
X$17143 \$16 \$10860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17144 \$16 \$8734 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17145 \$16 \$10529 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17147 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$17148 \$153 \$8734 \$11983 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$17149 \$16 \$11979 \$16 \$153 \$11824 VNB sky130_fd_sc_hd__clkbuf_2
X$17151 \$153 \$11781 \$11780 \$11947 \$11782 \$11803 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$17152 \$16 \$11915 \$16 \$153 \$11945 VNB sky130_fd_sc_hd__clkbuf_2
X$17153 \$153 \$7834 \$8340 \$12119 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17154 \$16 \$12017 \$16 \$153 \$11772 VNB sky130_fd_sc_hd__clkbuf_2
X$17156 \$153 \$11781 \$11782 \$12017 \$11780 \$11803 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$17157 \$153 \$10361 \$12120 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$17158 \$16 \$10361 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17159 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17160 \$153 \$8157 \$8340 \$11942 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17162 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17163 \$153 \$8283 \$8340 \$12179 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17164 \$16 \$11942 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17166 \$16 \$10392 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17167 \$153 \$12000 \$11809 \$10392 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17168 \$16 \$12179 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17169 \$16 \$12162 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17170 \$153 \$11809 \$12162 \$12077 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$17171 \$16 \$11824 \$16 \$153 \$11827 VNB sky130_fd_sc_hd__inv_1
X$17174 \$153 \$12000 \$10815 \$11827 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17175 \$16 \$11824 \$11504 \$12077 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$17177 \$16 \$11930 \$11504 \$12052 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$17178 \$16 \$11824 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17180 \$153 \$11629 \$11842 \$12052 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$17181 \$153 \$11703 \$10376 \$11515 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17182 \$153 \$11628 \$12009 \$11980 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$17184 \$16 \$11842 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17185 \$16 \$10392 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17186 \$153 \$11554 \$10560 \$11016 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17187 \$153 \$12001 \$11628 \$10617 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17188 \$153 \$12061 \$11628 \$10392 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17189 \$16 \$10739 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17191 \$153 \$12001 \$10560 \$11829 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17192 \$153 \$12122 \$11881 \$12121 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17193 \$153 \$12061 \$10815 \$11829 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17194 \$153 \$12145 \$11942 \$12121 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17195 \$16 \$12120 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17196 \$153 \$12123 \$12182 \$12121 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17198 \$153 \$11981 \$10815 \$11678 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17201 \$153 \$11916 \$10560 \$11678 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17202 \$16 \$12032 \$11504 \$12078 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$17203 \$153 \$11709 \$12198 \$12078 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$17204 \$16 \$11945 \$11504 \$12053 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$17206 \$153 \$11917 \$10376 \$11678 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17207 \$16 \$12120 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17208 \$153 \$12124 \$12087 \$12120 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17209 \$16 \$11945 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17211 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$17213 \$153 \$12035 \$12371 \$12147 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17214 \$16 \$12050 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17215 \$16 \$12220 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17216 \$153 \$12087 \$12050 \$12125 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$17217 \$153 \$11918 \$10587 \$11680 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17218 \$16 \$10736 \$12018 \$12146 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$17220 \$153 \$11920 \$10815 \$11680 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17221 \$16 \$12010 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17222 \$153 \$12126 \$12087 \$12010 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17223 \$153 \$12055 \$11681 \$10392 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17224 \$16 \$10981 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17225 \$16 \$10661 \$12018 \$12079 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$17226 \$16 \$10392 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17227 \$153 \$12088 \$10981 \$12079 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$17230 \$153 \$11982 \$10587 \$11730 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17232 \$16 \$12010 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17234 \$153 \$12080 \$12088 \$12010 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17236 \$153 \$12002 \$12088 \$11983 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17238 \$16 \$11983 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17239 \$153 \$11984 \$10560 \$11730 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17240 \$153 \$12080 \$11942 \$12127 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17241 \$153 \$12002 \$11881 \$12127 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17243 \$16 \$10853 \$12018 \$12128 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$17244 \$153 \$12036 \$12089 \$11983 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17245 \$153 \$12054 \$11881 \$12147 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17247 \$16 \$10853 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17249 \$153 \$12036 \$11881 \$11958 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17251 \$16 \$12010 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17252 \$16 \$12120 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17253 \$153 \$11957 \$12089 \$12010 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17254 \$153 \$11588 \$11776 \$11790 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$17255 \$16 \$11983 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17257 \$153 \$12037 \$10860 \$12062 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$17259 \$16 \$10529 \$12018 \$12062 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$17260 \$153 \$12129 \$12037 \$11983 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17261 \$153 \$12038 \$12339 \$11958 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17262 \$153 \$12039 \$12037 \$12010 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17263 \$16 \$12010 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17264 \$16 \$10860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17265 \$16 \$11390 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17267 \$16 \$10529 \$16 \$153 \$12011 VNB sky130_fd_sc_hd__inv_1
X$17268 \$16 \$10529 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17269 \$16 \$11390 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17270 \$153 \$12039 \$11942 \$12011 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17272 \$16 \$12384 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17273 \$153 \$12081 \$12037 \$12384 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17274 \$153 \$11392 \$10587 \$11390 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17275 \$16 \$11627 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17278 \$16 \$11390 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17279 \$153 \$11464 \$10815 \$11461 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17280 \$153 \$12081 \$12179 \$12011 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17281 \$153 \$11325 \$10376 \$11461 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17283 \$153 \$11388 \$10587 \$11461 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17284 \$153 \$10426 \$10815 \$10801 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17285 \$153 \$11175 \$10560 \$11461 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17287 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$17288 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$17289 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$17290 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$17291 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$17292 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$17293 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$17294 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$17295 \$153 \$9268 \$9458 \$8950 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17296 \$153 \$9062 \$9458 \$8715 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17297 \$153 \$8680 \$9458 \$9129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17298 \$16 \$8715 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17299 \$16 \$8950 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17300 \$16 \$8828 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17302 \$153 \$8896 \$9458 \$8828 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17303 \$16 \$8580 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17304 \$153 \$8979 \$9458 \$8724 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17305 \$153 \$9064 \$9458 \$9026 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17307 \$153 \$9065 \$9458 \$8436 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17308 \$153 \$9736 \$8209 \$9392 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17309 \$153 \$9545 \$8457 \$9392 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17310 \$16 \$7381 \$16 \$153 \$8679 VNB sky130_fd_sc_hd__inv_1
X$17311 \$153 \$9330 \$9469 \$9129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17312 \$16 \$9026 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17313 \$16 \$8436 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17314 \$16 \$8001 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17316 \$16 \$7884 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17317 \$16 \$7547 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17318 \$16 \$7381 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17319 \$153 \$9471 \$9469 \$8950 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17320 \$16 \$9129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17321 \$153 \$9470 \$8885 \$9270 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17323 \$153 \$9471 \$8912 \$9270 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17324 \$16 \$8950 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17325 \$153 \$9269 \$9469 \$8724 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17327 \$153 \$9469 \$8438 \$9472 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$17328 \$153 \$9473 \$9543 \$8724 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17329 \$153 \$9448 \$8457 \$9583 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17330 \$16 \$8003 \$9547 \$9472 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$17331 \$153 \$9473 \$8457 \$9449 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17333 \$16 \$8724 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17334 \$153 \$9546 \$8194 \$9449 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17335 \$153 \$9543 \$7655 \$9474 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$17336 \$16 \$7922 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17337 \$16 \$7655 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17338 \$153 \$9564 \$9543 \$9026 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17339 \$16 \$9220 \$16 \$153 \$9547 VNB sky130_fd_sc_hd__clkbuf_2
X$17342 \$153 \$9412 \$8737 \$9136 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17343 \$16 \$7922 \$16 \$153 \$9449 VNB sky130_fd_sc_hd__inv_1
X$17344 \$16 \$9026 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17345 \$16 \$7922 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17347 \$153 \$9508 \$9459 \$8950 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17348 \$153 \$9354 \$9459 \$9026 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17349 \$153 \$9475 \$9459 \$8828 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17350 \$16 \$9026 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17353 \$16 \$8436 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17355 \$16 \$8828 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17356 \$153 \$9413 \$9459 \$9129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17357 \$153 \$8910 \$8885 \$7816 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17358 \$16 \$7973 \$9260 \$9476 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$17360 \$16 \$7663 \$9260 \$9530 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$17362 \$153 \$9459 \$8117 \$9476 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$17363 \$153 \$9606 \$7887 \$9530 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$17364 \$16 \$9414 \$16 \$153 \$9200 VNB sky130_fd_sc_hd__clkbuf_2
X$17365 \$16 \$9414 \$16 \$153 \$3198 VNB sky130_fd_sc_hd__clkbuf_2
X$17368 \$153 \$9395 \$9334 \$8580 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17369 \$153 \$9509 \$8737 \$9322 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17372 \$16 \$8950 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17373 \$16 \$7887 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17374 \$16 \$8580 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17375 \$153 \$9509 \$9334 \$9129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17376 \$153 \$9565 \$9606 \$8724 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17377 \$16 \$7992 \$9260 \$9450 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$17378 \$16 \$7663 \$16 \$153 \$9585 VNB sky130_fd_sc_hd__inv_1
X$17380 \$153 \$9531 \$9334 \$8950 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17382 \$153 \$9334 \$8119 \$9450 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$17383 \$153 \$9460 \$8885 \$9322 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17384 \$153 \$9531 \$8912 \$9322 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17385 \$153 \$9415 \$8457 \$9322 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17386 \$16 \$8950 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17387 \$16 \$8125 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17389 \$16 \$7663 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17390 \$16 \$8715 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17392 \$153 \$9566 \$9384 \$8715 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17393 \$153 \$9477 \$9384 \$8580 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17394 \$16 \$8580 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17395 \$16 \$6887 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17396 \$16 \$8119 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17397 \$16 \$7535 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17398 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$17400 \$153 \$9532 \$9384 \$9026 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17402 \$153 \$9477 \$8194 \$9396 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17403 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$17404 \$16 \$9129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17405 \$153 \$9510 \$9384 \$8950 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17406 \$153 \$9532 \$8726 \$9396 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17407 \$16 \$9026 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17409 \$16 \$8950 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17412 \$153 \$9510 \$8912 \$9396 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17413 \$153 \$9398 \$9384 \$9129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17415 \$16 \$7922 \$9371 \$9568 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$17416 \$153 \$9416 \$8277 \$9417 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17418 \$153 \$9478 \$8727 \$9417 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17419 \$153 \$9478 \$9356 \$8886 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17421 \$153 \$9479 \$9356 \$8816 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17423 \$16 \$7922 \$16 \$153 \$9533 VNB sky130_fd_sc_hd__inv_1
X$17424 \$153 \$9479 \$8804 \$9417 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17425 \$153 \$9548 \$8727 \$9533 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17426 \$16 \$8816 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17427 \$16 \$8886 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17428 \$16 \$8890 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17430 \$16 \$7922 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17432 \$153 \$9549 \$8614 \$9417 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17433 \$153 \$9480 \$9356 \$8898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17434 \$16 \$8647 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17435 \$16 \$9569 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17436 \$16 \$8898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17437 \$153 \$9418 \$9356 \$8686 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17438 \$153 \$9480 \$8789 \$9417 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17440 \$153 \$9140 \$9356 \$8728 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17441 \$153 \$9534 \$8651 \$9451 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17443 \$153 \$9481 \$8438 \$9419 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$17444 \$153 \$9461 \$8818 \$9451 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17445 \$153 \$9482 \$9481 \$8556 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17447 \$153 \$9337 \$9481 \$8728 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17448 \$16 \$8556 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17449 \$153 \$9462 \$8804 \$9186 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17451 \$153 \$9483 \$9481 \$8647 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17452 \$16 \$8003 \$16 \$153 \$9186 VNB sky130_fd_sc_hd__inv_1
X$17455 \$16 \$8686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17456 \$153 \$9483 \$8614 \$9186 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17457 \$16 \$8647 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17458 \$16 \$9371 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17459 \$16 \$8297 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17460 \$153 \$9485 \$9484 \$8647 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17462 \$153 \$9399 \$9484 \$8890 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17463 \$16 \$8647 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17465 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$17466 \$16 \$8890 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17467 \$16 \$8144 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17468 \$16 \$8144 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17470 \$153 \$9511 \$9484 \$8686 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17471 \$153 \$9386 \$9484 \$8556 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17473 \$16 \$9273 \$16 \$153 \$9400 VNB sky130_fd_sc_hd__clkbuf_2
X$17474 \$153 \$9511 \$8651 \$9373 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17476 \$16 \$8686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17477 \$16 \$7973 \$9400 \$9486 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$17478 \$16 \$8556 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17479 \$153 \$9487 \$8117 \$9486 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$17480 \$153 \$9512 \$9487 \$8556 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17482 \$153 \$9464 \$9487 \$8686 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17483 \$16 \$9550 \$16 \$153 \$9273 VNB sky130_fd_sc_hd__clkbuf_2
X$17486 \$153 \$9513 \$9487 \$8728 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17487 \$153 \$9463 \$8119 \$9420 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$17488 \$16 \$9550 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17489 \$16 \$8686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17490 \$16 \$8728 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17492 \$153 \$9401 \$9463 \$8816 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17493 \$16 \$7973 \$16 \$153 \$9488 VNB sky130_fd_sc_hd__inv_1
X$17496 \$153 \$9514 \$9463 \$8898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17497 \$153 \$9514 \$8789 \$9421 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17498 \$153 \$9402 \$9463 \$8886 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17499 \$16 \$8898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17500 \$16 \$8816 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17501 \$16 \$8647 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17502 \$16 \$8556 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17504 \$153 \$9403 \$7887 \$9422 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$17505 \$153 \$9515 \$9463 \$8890 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17506 \$153 \$9570 \$9403 \$8647 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17508 \$16 \$7663 \$16 \$153 \$9452 VNB sky130_fd_sc_hd__inv_1
X$17509 \$16 \$8890 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17510 \$16 \$7663 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17512 \$16 \$6753 \$9400 \$9489 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$17513 \$16 \$8647 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17514 \$153 \$9571 \$9403 \$8686 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17515 \$153 \$9423 \$8610 \$9452 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17516 \$16 \$8556 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17518 \$16 \$8686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17519 \$153 \$9490 \$9424 \$8686 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17520 \$16 \$8686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17521 \$16 \$8886 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17522 \$16 \$6887 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17523 \$16 \$7535 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17526 \$153 \$9516 \$9424 \$8556 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17527 \$153 \$9464 \$8651 \$9488 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17529 \$153 \$9425 \$8804 \$9300 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17530 \$16 \$8556 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17532 \$16 \$8647 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17533 \$153 \$9572 \$9424 \$8647 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17534 \$16 \$6753 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17536 \$153 \$9491 \$9424 \$8728 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17537 \$153 \$9517 \$9424 \$8890 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17538 \$153 \$9426 \$8789 \$9300 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17539 \$16 \$8728 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17541 \$16 \$7490 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17543 \$16 \$9031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17544 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$17545 \$153 \$9079 \$9404 \$9031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17546 \$153 \$9213 \$9404 \$8936 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17547 \$153 \$9552 \$8727 \$9300 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17548 \$16 \$8936 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17549 \$16 \$8807 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17551 \$16 \$8126 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17553 \$16 \$9133 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17554 \$153 \$9517 \$8277 \$9300 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17555 \$16 \$9278 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17556 \$16 \$7347 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17557 \$153 \$8990 \$9404 \$9045 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17558 \$153 \$9722 \$8676 \$9453 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17559 \$153 \$9404 \$7852 \$9427 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$17560 \$16 \$9045 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17561 \$16 \$9188 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17563 \$16 \$7793 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17565 \$16 \$8078 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17566 \$16 \$7852 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17567 \$16 \$8819 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17568 \$16 \$9045 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17570 \$16 \$8936 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17571 \$153 \$9342 \$9405 \$9045 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17572 \$153 \$9343 \$9405 \$8936 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17573 \$153 \$9341 \$9405 \$8807 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17574 \$16 \$8187 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17577 \$153 \$9428 \$9047 \$9324 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17579 \$153 \$9492 \$9278 \$9324 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17580 \$16 \$9188 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17581 \$153 \$9492 \$9405 \$9275 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17582 \$153 \$9493 \$8900 \$9188 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17584 \$153 \$8916 \$9405 \$9188 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17586 \$153 \$9454 \$9133 \$9587 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17587 \$16 \$8361 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17588 \$153 \$9494 \$9081 \$8936 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17589 \$153 \$9494 \$8842 \$9276 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17591 \$16 \$8361 \$16 \$153 \$9455 VNB sky130_fd_sc_hd__clkbuf_2
X$17592 \$16 \$8936 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17593 \$153 \$9429 \$9252 \$9276 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17595 \$16 \$9455 \$16 \$153 \$9518 VNB sky130_fd_sc_hd__clkbuf_2
X$17596 \$153 \$9496 \$9081 \$9045 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17598 \$153 \$9495 \$9081 \$8807 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17601 \$153 \$9553 \$8676 \$9695 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17602 \$153 \$9496 \$9174 \$9276 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17604 \$153 \$9495 \$8676 \$9276 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17605 \$153 \$9554 \$9544 \$9045 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17606 \$16 \$9045 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17607 \$16 \$8807 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17608 \$16 \$9253 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17609 \$16 \$8044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17610 \$153 \$9554 \$9174 \$9465 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17612 \$153 \$9497 \$8676 \$9465 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17613 \$16 \$7904 \$16 \$153 \$9465 VNB sky130_fd_sc_hd__inv_1
X$17615 \$16 \$8807 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17616 \$16 \$7904 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17617 \$16 \$9045 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17618 \$153 \$9498 \$9466 \$8807 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17619 \$153 \$9432 \$9466 \$9045 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17621 \$16 \$9031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17622 \$153 \$9519 \$9466 \$9031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17623 \$153 \$9519 \$9133 \$9325 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17624 \$153 \$9573 \$9466 \$9275 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17625 \$153 \$9498 \$8676 \$9325 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17627 \$16 \$9455 \$16 \$153 \$9733 VNB sky130_fd_sc_hd__clkbuf_2
X$17630 \$16 \$7691 \$8960 \$9520 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$17632 \$16 \$8936 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17633 \$153 \$9574 \$9433 \$9188 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17634 \$153 \$9387 \$9433 \$8936 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17635 \$16 \$8772 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17636 \$16 \$9188 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17637 \$16 \$7691 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17639 \$16 \$9045 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17640 \$16 \$9031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17641 \$153 \$9522 \$9433 \$9045 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17643 \$153 \$9575 \$9433 \$9031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17644 \$16 \$7915 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17645 \$153 \$9522 \$9174 \$9521 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17646 \$16 \$8936 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17647 \$153 \$9361 \$8917 \$9033 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17649 \$16 \$9214 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17651 \$153 \$9523 \$9408 \$9214 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17652 \$153 \$9435 \$9408 \$8936 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17653 \$153 \$9523 \$9047 \$9409 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17654 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$17655 \$16 \$8265 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17656 \$16 \$9045 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17657 \$153 \$9499 \$9408 \$9045 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17659 \$16 \$8359 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17661 \$153 \$9434 \$8676 \$9409 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17663 \$16 \$8351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17664 \$153 \$9499 \$9174 \$9409 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17665 \$16 \$7695 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17666 \$153 \$9524 \$8351 \$9576 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$17667 \$16 \$9253 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17668 \$16 \$8101 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17670 \$16 \$9214 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17672 \$153 \$9500 \$9347 \$9214 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17673 \$153 \$9535 \$9524 \$9045 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17674 \$153 \$9535 \$9174 \$9555 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17675 \$153 \$9500 \$9047 \$9328 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17676 \$16 \$9031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17678 \$16 \$8936 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17679 \$153 \$9525 \$9347 \$9031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17681 \$153 \$9577 \$9524 \$8936 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17682 \$153 \$9309 \$8842 \$9328 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17683 \$153 \$9525 \$9133 \$9328 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17684 \$16 \$8359 \$16 \$153 \$9555 VNB sky130_fd_sc_hd__inv_1
X$17685 \$153 \$9556 \$8676 \$9555 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17688 \$16 \$7793 \$8824 \$9438 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$17689 \$16 \$7793 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17690 \$153 \$9578 \$9467 \$9134 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17691 \$153 \$9410 \$9467 \$8927 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17693 \$16 \$8927 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17694 \$153 \$9526 \$9467 \$9035 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17695 \$16 \$9134 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17698 \$16 \$8192 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17699 \$16 \$7386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17701 \$153 \$9526 \$8977 \$9439 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17703 \$153 \$9350 \$9467 \$9034 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17704 \$153 \$9579 \$9467 \$8844 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17706 \$16 \$9034 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17707 \$16 \$9154 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17709 \$16 \$7956 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17710 \$16 \$8844 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17711 \$16 \$7076 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17712 \$16 \$8429 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17713 \$153 \$9456 \$9256 \$9329 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17714 \$16 \$8429 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17715 \$153 \$9536 \$9122 \$9329 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17716 \$153 \$9501 \$9441 \$8844 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17717 \$153 \$9557 \$8996 \$9329 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17719 \$153 \$9536 \$9441 \$9134 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17720 \$153 \$9501 \$8965 \$9329 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17721 \$16 \$8844 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17722 \$16 \$8927 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17723 \$16 \$9035 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17725 \$16 \$9154 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17726 \$153 \$9502 \$9103 \$9329 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17727 \$153 \$9502 \$9441 \$9154 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17729 \$153 \$9503 \$9441 \$9035 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17730 \$153 \$9558 \$8996 \$9560 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17731 \$153 \$9559 \$9122 \$9560 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17732 \$153 \$9503 \$8977 \$9329 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17733 \$153 \$9468 \$8250 \$9457 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$17734 \$16 \$8136 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17738 \$153 \$9561 \$9059 \$9560 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17740 \$16 \$8044 \$9675 \$9457 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$17741 \$16 \$8927 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17742 \$153 \$9504 \$9468 \$8927 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17743 \$16 \$8250 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17745 \$153 \$9504 \$9256 \$9411 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17747 \$16 \$8844 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17748 \$153 \$9537 \$9468 \$9134 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17749 \$16 \$9134 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17751 \$16 \$9035 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17752 \$153 \$9389 \$9468 \$9035 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17753 \$153 \$9537 \$9122 \$9411 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17754 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$17755 \$16 \$9034 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17756 \$16 \$8844 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17758 \$153 \$9505 \$9468 \$8844 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17759 \$153 \$9538 \$9468 \$9034 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17760 \$153 \$9538 \$9059 \$9411 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17761 \$153 \$9505 \$8965 \$9411 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17762 \$16 \$9191 \$16 \$153 \$9562 VNB sky130_fd_sc_hd__clkbuf_2
X$17763 \$16 \$8927 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17765 \$16 \$8844 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17767 \$153 \$9527 \$9364 \$8927 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17768 \$153 \$9539 \$9364 \$8844 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17770 \$153 \$9365 \$9059 \$9280 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17771 \$153 \$9539 \$8965 \$9280 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17772 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$17774 \$153 \$9563 \$9103 \$9280 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17775 \$153 \$9443 \$8996 \$9280 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17776 \$16 \$9154 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17777 \$153 \$9506 \$9316 \$9154 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17779 \$16 \$9035 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17780 \$153 \$9507 \$9316 \$9035 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17782 \$153 \$9507 \$8977 \$9239 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17783 \$16 \$8316 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17784 \$16 \$9134 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17785 \$16 \$8893 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17786 \$153 \$9540 \$9316 \$8893 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17787 \$153 \$9506 \$9103 \$9239 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17788 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$17789 \$153 \$9444 \$9059 \$9239 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17790 \$16 \$8266 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17791 \$16 \$8351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17793 \$153 \$9581 \$8351 \$9580 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$17794 \$16 \$8101 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17795 \$16 \$7695 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17797 \$16 \$8893 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17798 \$153 \$9445 \$9391 \$8893 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17799 \$16 \$8879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17800 \$153 \$9541 \$9391 \$8879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17802 \$16 \$8265 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17803 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$17805 \$153 \$9541 \$8923 \$9366 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17806 \$16 \$8927 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17807 \$153 \$9528 \$9391 \$8927 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17808 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$17810 \$153 \$9542 \$8965 \$9366 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17811 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$17812 \$16 \$9035 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17814 \$153 \$9529 \$9391 \$9035 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17816 \$16 \$8844 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17817 \$153 \$9542 \$9391 \$8844 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17818 \$16 \$9154 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17819 \$153 \$9367 \$8965 \$9192 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17820 \$153 \$9529 \$8977 \$9366 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17822 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$17823 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$17825 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$17826 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$17827 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$17828 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$17830 \$153 \$10328 \$10327 \$10006 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17831 \$153 \$10255 \$10276 \$10006 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17832 \$153 \$10301 \$10256 \$10295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17833 \$153 \$10225 \$10256 \$10368 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17835 \$153 \$10225 \$10303 \$10245 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17837 \$153 \$10301 \$10276 \$10245 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17838 \$16 \$10368 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17839 \$16 \$10295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17840 \$153 \$10208 \$10256 \$10200 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17842 \$153 \$10329 \$10318 \$10245 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17843 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$17844 \$16 \$10200 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17848 \$153 \$10271 \$10256 \$10226 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17849 \$153 \$10271 \$10161 \$10245 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17850 \$153 \$10347 \$10276 \$10210 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17851 \$16 \$10226 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17853 \$153 \$10209 \$10250 \$10368 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17854 \$153 \$10272 \$10161 \$10210 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17856 \$16 \$10348 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17857 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$17858 \$153 \$10302 \$10330 \$10210 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17859 \$153 \$10272 \$10250 \$10226 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17860 \$153 \$10087 \$10250 \$10200 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17861 \$16 \$10368 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17862 \$16 \$10226 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17865 \$153 \$10257 \$10318 \$10210 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17866 \$16 \$10646 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17867 \$16 \$10200 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17869 \$16 \$10539 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17871 \$153 \$10227 \$10251 \$10226 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17872 \$153 \$10296 \$10251 \$10295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17873 \$153 \$10258 \$10318 \$10211 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17874 \$16 \$10295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17876 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$17877 \$153 \$10136 \$10251 \$10200 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17878 \$16 \$10226 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17880 \$153 \$10273 \$10251 \$10368 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17881 \$16 \$10200 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17883 \$153 \$10273 \$10303 \$10211 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17884 \$16 \$10368 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17886 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$17889 \$153 \$10349 \$10259 \$10226 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17890 \$153 \$10274 \$10259 \$10368 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17891 \$16 \$10368 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17892 \$16 \$10226 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17893 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$17895 \$16 \$9026 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17896 \$153 \$10228 \$10259 \$10200 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17899 \$153 \$10274 \$10303 \$10246 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17900 \$153 \$10349 \$10161 \$10246 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17901 \$153 \$10228 \$10088 \$10246 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17902 \$16 \$10200 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17903 \$16 \$6057 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17904 \$16 \$6057 \$16 \$153 \$8361 VNB sky130_fd_sc_hd__clkbuf_2
X$17906 \$153 \$10187 \$10199 \$10226 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17909 \$153 \$10213 \$10199 \$10368 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17910 \$153 \$10304 \$10199 \$10295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17912 \$153 \$6693 \$8838 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$17914 \$153 \$10186 \$10088 \$10212 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17915 \$16 \$10143 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17916 \$153 \$10304 \$10276 \$10212 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17918 \$153 \$10275 \$10252 \$10295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17920 \$153 \$10305 \$10252 \$10200 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17922 \$153 \$10229 \$10252 \$10226 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17924 \$153 \$10305 \$10088 \$10331 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17925 \$153 \$10229 \$10161 \$10331 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17926 \$153 \$10275 \$10276 \$10331 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17927 \$153 \$8839 \$10226 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$17928 \$16 \$8839 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17931 \$153 \$10332 \$10303 \$10331 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17932 \$153 \$10333 \$10318 \$10331 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17933 \$153 \$9802 \$8457 \$9866 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17934 \$16 \$8436 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17935 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$17936 \$16 \$6722 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17937 \$153 \$9339 \$10368 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$17939 \$153 \$10042 \$10200 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$17940 \$16 \$9339 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17941 \$153 \$10351 \$10276 \$10334 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17942 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17943 \$16 \$10042 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17945 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17946 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17948 \$153 \$10306 \$8340 \$10318 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17949 \$153 \$10079 \$8340 \$10303 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17950 \$153 \$10036 \$4037 \$10230 \$10306 \$10319 \$8956 \$10007 \$16 \$16
+ VNB sky130_fd_sc_hd__mux4_1
X$17951 \$153 \$9685 \$8457 \$9567 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17952 \$16 \$10303 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17954 \$16 \$10161 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17955 \$16 \$8726 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17957 \$16 \$10276 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17958 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17959 \$16 \$8956 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17960 \$153 \$10018 \$8340 \$10276 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17961 \$153 \$10036 \$4039 \$10119 \$10433 \$10260 \$8788 \$10007 \$16 \$16
+ VNB sky130_fd_sc_hd__mux4_1
X$17962 \$16 \$10606 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17966 \$16 \$6649 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17967 \$153 \$10297 \$9900 \$8890 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17968 \$153 \$6649 \$9747 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$17969 \$153 \$10353 \$10320 \$10298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17970 \$16 \$8890 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17971 \$16 \$8114 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17973 \$16 \$8788 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17974 \$16 \$8955 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17976 \$153 \$10162 \$8804 \$9868 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17977 \$153 \$10335 \$10098 \$10369 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17978 \$153 \$6799 \$9138 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$17979 \$153 \$10297 \$8277 \$9868 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17980 \$16 \$10382 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17984 \$153 \$10336 \$10098 \$10337 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$17985 \$153 \$10214 \$9794 \$8890 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17987 \$153 \$10307 \$10400 \$10470 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17988 \$16 \$6799 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17989 \$16 \$8890 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17992 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$17993 \$16 \$10298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17994 \$16 \$10470 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17995 \$153 \$10137 \$9795 \$8890 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$17997 \$153 \$6669 \$8301 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$17998 \$16 \$8890 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$17999 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$18000 \$153 \$10163 \$8804 \$9720 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18002 \$153 \$10355 \$10309 \$10339 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18004 \$153 \$10150 \$9796 \$8816 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18005 \$153 \$10308 \$10380 \$10298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18006 \$16 \$8816 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18007 \$153 \$10308 \$10401 \$10339 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18011 \$153 \$6653 \$8670 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$18012 \$16 \$10298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18013 \$153 \$10310 \$9811 \$8890 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18014 \$16 \$6653 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18016 \$16 \$10338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18017 \$153 \$10164 \$8804 \$9586 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18018 \$16 \$10321 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18020 \$153 \$10356 \$10309 \$10515 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18022 \$153 \$10167 \$3240 \$8760 \$10215 \$9886 \$10081 \$10082 \$16 \$16
+ VNB sky130_fd_sc_hd__mux4_1
X$18023 \$153 \$10167 \$3646 \$8607 \$10321 \$10322 \$10299 \$10082 \$16 \$16
+ VNB sky130_fd_sc_hd__mux4_1
X$18025 \$153 \$10167 \$3842 \$8411 \$10165 \$10253 \$9970 \$10082 \$16 \$16
+ VNB sky130_fd_sc_hd__mux4_1
X$18027 \$16 \$6654 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18028 \$153 \$6654 \$8516 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$18029 \$153 \$10248 \$10247 \$10249 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18031 \$16 \$10261 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18033 \$16 \$10357 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18035 \$153 \$10341 \$10098 \$10249 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18036 \$153 \$10167 \$4340 \$8555 \$10261 \$10262 \$10153 \$10082 \$16 \$16
+ VNB sky130_fd_sc_hd__mux4_1
X$18037 \$153 \$10342 \$10323 \$10338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18038 \$16 \$8487 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18039 \$16 \$6735 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18042 \$153 \$6735 \$8364 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$18043 \$153 \$10358 \$10323 \$10298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18044 \$153 \$10342 \$10309 \$10343 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18045 \$153 \$10097 \$10298 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$18047 \$16 \$9997 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18049 \$153 \$9997 \$10382 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$18050 \$153 \$9848 \$8727 \$9746 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18051 \$16 \$10097 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18052 \$153 \$10527 \$8890 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$18054 \$16 \$10408 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18055 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18057 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18058 \$153 \$10254 \$8340 \$8727 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18059 \$153 \$10264 \$8340 \$10344 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18060 \$153 \$10042 \$10473 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$18062 \$153 \$9998 \$8727 \$9845 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18063 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18064 \$153 \$10277 \$8340 \$8277 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18065 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18067 \$153 \$10061 \$8340 \$10309 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18068 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18070 \$153 \$9971 \$9252 \$9453 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18071 \$153 \$10101 \$8340 \$10247 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18072 \$153 \$10299 \$8340 \$9047 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18073 \$153 \$10046 \$8842 \$9453 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18074 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18078 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18079 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18080 \$153 \$10278 \$8340 \$8789 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18082 \$153 \$10263 \$10021 \$9275 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18083 \$153 \$10263 \$9278 \$10216 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18084 \$16 \$10309 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18085 \$16 \$10344 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18086 \$16 \$10516 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18087 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18089 \$153 \$10359 \$10021 \$9188 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18091 \$153 \$10279 \$10021 \$9253 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18092 \$153 \$10279 \$9252 \$10216 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18093 \$16 \$9253 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18095 \$16 \$9214 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18096 \$153 \$10280 \$10000 \$9214 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18097 \$16 \$9252 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18098 \$16 \$8673 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18100 \$153 \$10359 \$8917 \$10216 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18102 \$16 \$6911 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18103 \$16 \$9253 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18105 \$153 \$10281 \$10000 \$9253 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18106 \$153 \$10217 \$10000 \$9275 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18108 \$16 \$8313 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18109 \$16 \$9275 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18112 \$16 \$9188 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18113 \$16 \$9214 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18114 \$153 \$10218 \$10083 \$9214 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18115 \$153 \$10360 \$10083 \$9188 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18116 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$18117 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$18118 \$16 \$7996 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18119 \$16 \$9253 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18120 \$16 \$9275 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18122 \$153 \$10312 \$10083 \$9253 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18123 \$153 \$10232 \$10083 \$9275 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18124 \$153 \$10312 \$9252 \$9953 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18125 \$153 \$10232 \$9278 \$9953 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18126 \$16 \$9275 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18128 \$153 \$10313 \$9934 \$9253 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18130 \$153 \$10233 \$9934 \$9275 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18131 \$153 \$10313 \$9252 \$9927 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18132 \$153 \$10233 \$9278 \$9927 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18133 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$18135 \$16 \$9188 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18136 \$16 \$9275 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18138 \$153 \$10234 \$10022 \$9275 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18139 \$153 \$10314 \$10022 \$9188 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18140 \$153 \$10234 \$9278 \$10009 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18141 \$153 \$10071 \$8676 \$10009 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18142 \$16 \$9214 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18143 \$153 \$7089 \$8416 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$18145 \$153 \$10156 \$10022 \$9214 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18146 \$153 \$10282 \$10024 \$9253 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18147 \$16 \$7089 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18148 \$153 \$10235 \$8917 \$10104 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18150 \$153 \$10282 \$9252 \$10104 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18151 \$153 \$10283 \$10024 \$9214 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18152 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$18154 \$153 \$10283 \$9047 \$10104 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18155 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$18156 \$16 \$7075 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18157 \$153 \$10125 \$9133 \$10104 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18159 \$153 \$7075 \$8734 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$18160 \$153 \$10219 \$10157 \$9253 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18161 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$18162 \$16 \$9253 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18164 \$16 \$9214 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18165 \$16 \$9275 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18167 \$153 \$10284 \$10157 \$9275 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18168 \$153 \$10196 \$10157 \$9214 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18169 \$153 \$10284 \$9278 \$9872 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18171 \$16 \$10300 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18172 \$16 \$9253 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18173 \$16 \$9214 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18174 \$153 \$10237 \$10010 \$9214 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18176 \$16 \$9031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18178 \$153 \$10236 \$10010 \$9253 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18179 \$153 \$10315 \$10388 \$10300 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18180 \$16 \$10192 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18181 \$153 \$10221 \$10010 \$9275 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18185 \$153 \$10075 \$3248 \$10278 \$10384 \$10316 \$10324 \$10220 \$16 \$16
+ VNB sky130_fd_sc_hd__mux4_1
X$18186 \$153 \$10075 \$3964 \$10192 \$10265 \$10266 \$10174 \$10220 \$16 \$16
+ VNB sky130_fd_sc_hd__mux4_1
X$18187 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18188 \$153 \$10267 \$8340 \$9059 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18191 \$153 \$10075 \$3087 \$10254 \$10264 \$10268 \$10267 \$10220 \$16 \$16
+ VNB sky130_fd_sc_hd__mux4_1
X$18192 \$153 \$10324 \$8340 \$8977 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18193 \$16 \$10264 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18194 \$16 \$10254 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18195 \$16 \$9059 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18196 \$16 \$10285 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18198 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$18199 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18200 \$16 \$8977 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18201 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$18203 \$153 \$7094 \$10238 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$18204 \$153 \$10408 \$9035 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$18205 \$16 \$7094 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18207 \$153 \$10286 \$9913 \$9134 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18208 \$153 \$10527 \$9134 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$18209 \$16 \$9134 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18210 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$18211 \$16 \$10527 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18212 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$18214 \$153 \$10205 \$9034 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$18216 \$153 \$7179 \$10205 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$18217 \$153 \$10239 \$8923 \$10108 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18218 \$153 \$9983 \$9256 \$10108 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18220 \$153 \$10287 \$9940 \$9034 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18221 \$16 \$7179 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18222 \$16 \$10043 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18223 \$16 \$9034 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18225 \$153 \$10287 \$9059 \$10108 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18226 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$18227 \$153 \$10129 \$9122 \$10108 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18228 \$16 \$9034 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18229 \$153 \$10288 \$10025 \$9034 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18232 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$18233 \$153 \$7099 \$10097 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$18235 \$16 \$9134 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18236 \$153 \$10289 \$10025 \$9134 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18238 \$153 \$10097 \$10346 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$18239 \$16 \$7099 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18241 \$153 \$10097 \$8879 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$18242 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$18243 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$18244 \$16 \$9134 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18245 \$16 \$9034 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18247 \$153 \$10317 \$10085 \$9134 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18248 \$153 \$10241 \$10085 \$9034 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18249 \$153 \$10241 \$9059 \$10110 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18250 \$153 \$10317 \$9122 \$10110 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18251 \$16 \$9034 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18252 \$16 \$10222 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18255 \$153 \$10290 \$10111 \$9034 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18256 \$16 \$10326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18257 \$153 \$10363 \$10395 \$10326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18258 \$16 \$9035 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18259 \$153 \$10223 \$10111 \$9035 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18260 \$153 \$10242 \$8923 \$9988 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18263 \$153 \$10364 \$10325 \$10326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18264 \$153 \$10243 \$9122 \$9988 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18266 \$16 \$9035 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18267 \$16 \$10326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18268 \$153 \$10269 \$9122 \$9961 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18270 \$16 \$9134 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18271 \$153 \$10269 \$9860 \$9134 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18273 \$153 \$10291 \$9860 \$9035 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18275 \$153 \$10291 \$8977 \$9961 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18276 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$18277 \$16 \$9035 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18279 \$153 \$10224 \$10028 \$9035 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18280 \$16 \$8085 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18281 \$16 \$10346 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18282 \$16 \$8879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18284 \$153 \$10365 \$10028 \$8879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18285 \$16 \$9134 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18286 \$153 \$10292 \$10028 \$9134 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18287 \$153 \$10366 \$10028 \$9034 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18289 \$153 \$10270 \$9122 \$10005 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18290 \$16 \$10326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18291 \$16 \$9134 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18292 \$153 \$10270 \$9991 \$9134 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18293 \$153 \$10293 \$9991 \$8879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18294 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$18295 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$18297 \$153 \$10293 \$8923 \$10005 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18298 \$16 \$9034 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18299 \$153 \$10294 \$9991 \$9034 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18301 \$153 \$10294 \$9059 \$10005 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18302 \$153 \$10244 \$8977 \$10005 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18303 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$18306 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$18307 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$18308 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$18309 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$18310 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$18311 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$18314 \$153 \$8202 \$8113 \$6783 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18315 \$153 \$8201 \$8113 \$6981 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18317 \$153 \$8360 \$6930 \$8384 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18318 \$153 \$8292 \$8113 \$6784 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18320 \$16 \$6981 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18322 \$153 \$8292 \$6794 \$8034 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18323 \$16 \$6783 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18324 \$16 \$6784 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18325 \$153 \$8203 \$8113 \$6792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18326 \$153 \$8332 \$8331 \$6979 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18328 \$153 \$8113 \$8193 \$8270 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$18329 \$153 \$8332 \$6995 \$8384 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18330 \$16 \$8114 \$16 \$153 \$8034 VNB sky130_fd_sc_hd__inv_1
X$18331 \$153 \$8204 \$8333 \$6979 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18332 \$16 \$6792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18334 \$153 \$8293 \$8333 \$6792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18336 \$16 \$6979 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18337 \$16 \$6860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18338 \$16 \$8114 \$8024 \$8270 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$18339 \$153 \$8293 \$6719 \$8206 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18340 \$16 \$6792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18341 \$153 \$8294 \$8333 \$6783 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18343 \$153 \$8205 \$8333 \$6981 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18345 \$153 \$8294 \$6749 \$8206 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18346 \$16 \$8423 \$16 \$153 \$8206 VNB sky130_fd_sc_hd__inv_1
X$18347 \$16 \$6783 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18348 \$16 \$6981 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18350 \$153 \$8295 \$8115 \$6907 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18351 \$153 \$8385 \$8115 \$6860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18352 \$153 \$8228 \$6995 \$8036 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18353 \$16 \$6860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18355 \$16 \$8503 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18357 \$16 \$8271 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18358 \$153 \$8334 \$8115 \$6784 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18359 \$16 \$6907 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18361 \$16 \$8271 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18362 \$16 \$8271 \$16 \$153 \$8036 VNB sky130_fd_sc_hd__inv_1
X$18363 \$153 \$8141 \$6749 \$8036 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18364 \$153 \$8334 \$6794 \$8036 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18365 \$16 \$8144 \$8024 \$8229 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$18367 \$16 \$6784 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18370 \$153 \$8296 \$8230 \$6783 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18371 \$153 \$8336 \$8230 \$6860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18372 \$153 \$8296 \$6749 \$8208 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18373 \$16 \$6783 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18375 \$16 \$8144 \$16 \$153 \$8208 VNB sky130_fd_sc_hd__inv_1
X$18376 \$153 \$8298 \$8230 \$6981 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18378 \$153 \$8175 \$8230 \$6979 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18379 \$153 \$8298 \$6930 \$8208 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18380 \$16 \$6981 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18381 \$16 \$8361 \$16 \$153 \$7467 VNB sky130_fd_sc_hd__clkbuf_2
X$18382 \$16 \$7467 \$16 \$153 \$8195 VNB sky130_fd_sc_hd__clkbuf_2
X$18383 \$153 \$8337 \$8272 \$6783 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18384 \$16 \$6981 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18386 \$153 \$8757 \$8457 \$7816 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18387 \$153 \$8299 \$8272 \$6979 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18388 \$153 \$8337 \$6749 \$8363 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18389 \$153 \$8362 \$6930 \$8363 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18390 \$153 \$8300 \$8272 \$6792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18392 \$153 \$8299 \$6995 \$8363 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18394 \$153 \$8300 \$6719 \$8363 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18395 \$153 \$8272 \$8119 \$8273 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$18396 \$16 \$7992 \$8195 \$8273 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$18397 \$153 \$8210 \$8274 \$6792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18400 \$153 \$8231 \$8274 \$6783 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18401 \$16 \$6783 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18402 \$153 \$8274 \$8169 \$8168 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$18403 \$153 \$8231 \$6749 \$8196 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18404 \$153 \$8232 \$8274 \$6981 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18406 \$153 \$8178 \$8274 \$6979 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18407 \$153 \$8232 \$6930 \$8196 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18409 \$16 \$8121 \$7399 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$18410 \$153 \$8364 \$6979 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$18411 \$16 \$8120 \$16 \$153 \$7992 VNB sky130_fd_sc_hd__clkbuf_2
X$18412 \$16 \$8301 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18414 \$16 \$8064 \$16 \$153 \$7973 VNB sky130_fd_sc_hd__clkbuf_2
X$18415 \$16 \$8233 \$16 \$153 \$8118 VNB sky130_fd_sc_hd__clkbuf_2
X$18416 \$16 \$7944 \$16 \$153 \$8005 VNB sky130_fd_sc_hd__clkbuf_2
X$18417 \$16 \$8275 \$16 \$153 \$8121 VNB sky130_fd_sc_hd__clkbuf_2
X$18418 \$16 \$7786 \$16 \$153 \$7989 VNB sky130_fd_sc_hd__clkbuf_2
X$18419 \$16 \$8275 \$16 \$153 \$7945 VNB sky130_fd_sc_hd__clkbuf_2
X$18420 \$16 \$8065 \$16 \$153 \$8177 VNB sky130_fd_sc_hd__clkbuf_2
X$18421 \$16 \$8142 \$16 \$153 \$6753 VNB sky130_fd_sc_hd__clkbuf_2
X$18422 \$16 \$7889 \$16 \$153 \$8026 VNB sky130_fd_sc_hd__clkbuf_2
X$18423 \$16 \$8121 \$7335 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$18424 \$16 \$8143 \$16 \$153 \$7535 VNB sky130_fd_sc_hd__clkbuf_2
X$18425 \$16 \$8255 \$16 \$153 \$8271 VNB sky130_fd_sc_hd__clkbuf_2
X$18428 \$16 \$8234 \$16 \$153 \$8139 VNB sky130_fd_sc_hd__clkbuf_2
X$18429 \$16 \$8276 \$16 \$153 \$8114 VNB sky130_fd_sc_hd__clkbuf_2
X$18430 \$153 \$8276 \$8038 \$7990 \$8066 \$8067 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$18431 \$153 \$8234 \$8038 \$8066 \$8067 \$7990 \$16 \$16 VNB
+ sky130_fd_sc_hd__nor4b_2
X$18432 \$153 \$8038 \$8067 \$8255 \$8066 \$7990 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$18433 \$153 \$8066 \$8038 \$8106 \$8067 \$7990 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$18434 \$16 \$8114 \$7968 \$8386 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$18436 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18437 \$153 \$8366 \$8818 \$8256 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18438 \$153 \$8257 \$8277 \$8256 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18439 \$153 \$8213 \$8356 \$6862 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18440 \$153 \$8302 \$8356 \$6991 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18441 \$16 \$6991 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18442 \$153 \$8302 \$6992 \$8214 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18444 \$153 \$8367 \$6906 \$8214 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18445 \$16 \$7945 \$8025 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$18446 \$16 \$8114 \$16 \$153 \$8214 VNB sky130_fd_sc_hd__inv_1
X$18448 \$153 \$8303 \$8356 \$7060 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18449 \$16 \$6862 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18450 \$153 \$8258 \$8356 \$6771 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18452 \$153 \$8258 \$6865 \$8214 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18453 \$153 \$8303 \$6324 \$8214 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18454 \$16 \$7060 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18456 \$16 \$6771 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18457 \$153 \$8304 \$8147 \$7060 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18458 \$16 \$8139 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18459 \$16 \$8193 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18460 \$16 \$8114 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18461 \$153 \$8304 \$6324 \$8107 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18463 \$16 \$7060 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18464 \$153 \$8368 \$6867 \$8107 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18465 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$18466 \$153 \$8305 \$8147 \$6862 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18468 \$153 \$8369 \$7006 \$8107 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18469 \$153 \$8370 \$6865 \$8107 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18470 \$16 \$6862 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18471 \$16 \$8271 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18473 \$16 \$8297 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18474 \$16 \$6771 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18475 \$153 \$7707 \$8297 \$8235 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$18476 \$16 \$8335 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18477 \$153 \$8388 \$7947 \$6916 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18478 \$16 \$8423 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18480 \$16 \$8144 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18481 \$16 \$8271 \$16 \$153 \$8040 VNB sky130_fd_sc_hd__inv_1
X$18482 \$16 \$7521 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18484 \$153 \$8306 \$7947 \$6771 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18485 \$16 \$6916 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18486 \$16 \$8271 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18488 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$18489 \$16 \$7060 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18490 \$153 \$8306 \$6865 \$8040 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18491 \$153 \$8215 \$8278 \$6862 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18493 \$153 \$8505 \$8278 \$6754 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18495 \$16 \$6862 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18497 \$16 \$7466 \$8357 \$8307 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$18498 \$16 \$6754 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18499 \$153 \$8259 \$8278 \$6797 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18500 \$153 \$8216 \$8278 \$6991 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18501 \$153 \$8259 \$6906 \$8217 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18502 \$16 \$6991 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18505 \$16 \$8117 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18506 \$16 \$7973 \$16 \$153 \$8218 VNB sky130_fd_sc_hd__inv_1
X$18507 \$16 \$6797 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18508 \$153 \$8338 \$8279 \$7044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18510 \$153 \$8236 \$8279 \$6916 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18511 \$153 \$8371 \$6865 \$8218 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18512 \$16 \$6916 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18513 \$16 \$8119 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18515 \$16 \$8025 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18516 \$153 \$8339 \$8279 \$6862 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18517 \$153 \$8308 \$8279 \$6991 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18518 \$153 \$8308 \$6992 \$8218 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18519 \$16 \$6991 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18520 \$16 \$6862 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18521 \$153 \$8309 \$8025 \$8091 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$18524 \$16 \$6935 \$8357 \$8389 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$18526 \$153 \$8170 \$8309 \$6862 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18528 \$153 \$8310 \$8309 \$6797 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18529 \$153 \$8310 \$6906 \$8260 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18530 \$16 \$8125 \$16 \$153 \$7933 VNB sky130_fd_sc_hd__inv_1
X$18532 \$16 \$8118 \$16 \$153 \$8260 VNB sky130_fd_sc_hd__inv_1
X$18533 \$16 \$6797 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18534 \$16 \$6862 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18535 \$16 \$8125 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18536 \$16 \$6935 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18537 \$153 \$8237 \$8309 \$6754 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18538 \$16 \$8118 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18539 \$153 \$8390 \$8309 \$6991 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18540 \$153 \$8237 \$6756 \$8260 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18541 \$16 \$6991 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18544 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$18545 \$16 \$6754 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18546 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$18547 \$153 \$8311 \$8027 \$7044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18548 \$153 \$8320 \$6754 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$18549 \$16 \$7044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18552 \$16 \$8320 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18553 \$153 \$10311 \$6991 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$18555 \$153 \$8391 \$6862 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$18556 \$16 \$10311 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18557 \$16 \$8391 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18558 \$153 \$153 \$7490 \$8219 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18559 \$16 \$8347 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18560 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18562 \$153 \$153 \$7215 \$8219 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18563 \$153 \$153 \$7065 \$8219 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18564 \$153 \$8341 \$8340 \$7003 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18565 \$153 \$153 \$6582 \$8219 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18566 \$16 \$8078 \$16 \$153 \$8219 VNB sky130_fd_sc_hd__clkbuf_2
X$18567 \$16 \$7934 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18568 \$16 \$7239 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18569 \$16 \$6992 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18571 \$153 \$8312 \$8028 \$7239 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18572 \$153 \$8392 \$8028 \$7067 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18573 \$153 \$8127 \$8028 \$7029 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18574 \$153 \$8238 \$7327 \$7860 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18575 \$16 \$7067 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18577 \$153 \$8312 \$7482 \$7860 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18579 \$16 \$8187 \$16 \$153 \$7860 VNB sky130_fd_sc_hd__inv_1
X$18581 \$153 \$8128 \$7874 \$7067 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18582 \$16 \$8187 \$8280 \$8348 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$18583 \$153 \$8028 \$7839 \$8348 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$18584 \$16 \$7067 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18587 \$16 \$8187 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18588 \$16 \$7839 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18589 \$16 \$7386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18591 \$16 \$8220 \$8280 \$8261 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$18592 \$16 \$8220 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18593 \$153 \$8372 \$7327 \$8373 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18594 \$153 \$7874 \$9150 \$8261 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$18595 \$16 \$7029 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18596 \$16 \$7328 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18597 \$153 \$8374 \$7066 \$8373 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18598 \$16 \$8220 \$16 \$153 \$7924 VNB sky130_fd_sc_hd__inv_1
X$18599 \$153 \$8239 \$8183 \$7328 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18601 \$153 \$8130 \$8183 \$7082 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18602 \$153 \$8239 \$7366 \$8043 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18603 \$153 \$8375 \$7327 \$8043 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18604 \$16 \$8313 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18605 \$16 \$8044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18606 \$16 \$7067 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18607 \$16 \$7082 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18609 \$16 \$8313 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18610 \$153 \$8221 \$8183 \$7067 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18611 \$16 \$8393 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18612 \$16 \$7387 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18613 \$153 \$8394 \$8183 \$7387 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18614 \$16 \$8506 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18615 \$16 \$8044 \$8280 \$8262 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$18616 \$16 \$7996 \$8280 \$8395 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$18617 \$153 \$7876 \$8250 \$8262 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$18618 \$16 \$8730 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18621 \$16 \$7387 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18622 \$16 \$7904 \$8280 \$8240 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$18623 \$153 \$8314 \$8281 \$7082 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18624 \$153 \$8342 \$8281 \$7387 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18627 \$153 \$8342 \$7490 \$8263 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18628 \$16 \$7082 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18630 \$153 \$8282 \$7066 \$8263 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18631 \$153 \$8314 \$7065 \$8263 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18632 \$153 \$8223 \$8029 \$7082 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18633 \$16 \$7994 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18635 \$153 \$8376 \$7482 \$8222 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18636 \$16 \$8283 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18640 \$16 \$7328 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18641 \$153 \$8396 \$8029 \$7067 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18642 \$153 \$8284 \$7366 \$8222 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18643 \$153 \$8315 \$8184 \$7328 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18644 \$153 \$8241 \$7215 \$8047 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18645 \$153 \$8315 \$7366 \$8047 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18648 \$16 \$8285 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18649 \$16 \$8316 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18651 \$16 \$8316 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18652 \$153 \$8349 \$6582 \$8047 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18653 \$153 \$7203 \$7066 \$6656 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18654 \$153 \$8350 \$7482 \$8047 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18655 \$153 \$8242 \$7327 \$8047 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18656 \$16 \$6656 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18657 \$16 \$6656 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18658 \$16 \$7328 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18659 \$153 \$8286 \$7215 \$8264 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18661 \$153 \$8397 \$8030 \$7328 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18662 \$153 \$8243 \$7066 \$8264 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18663 \$153 \$8397 \$7366 \$8264 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18664 \$153 \$8160 \$6582 \$8264 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18666 \$153 \$8343 \$8358 \$7082 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18670 \$16 \$7387 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18671 \$153 \$8317 \$8030 \$7387 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18672 \$153 \$8343 \$7065 \$8527 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18674 \$16 \$8359 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18675 \$16 \$7239 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18676 \$16 \$7082 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18677 \$16 \$8265 \$16 \$153 \$8264 VNB sky130_fd_sc_hd__inv_1
X$18679 \$16 \$8351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18680 \$153 \$8131 \$8030 \$7239 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18682 \$153 \$8317 \$7490 \$8264 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18683 \$16 \$8359 \$8573 \$8352 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$18684 \$153 \$8244 \$7327 \$8264 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18685 \$153 \$7953 \$8351 \$8352 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$18687 \$16 \$8359 \$16 \$153 \$8048 VNB sky130_fd_sc_hd__inv_1
X$18690 \$16 \$8265 \$8573 \$8398 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$18691 \$16 \$8224 \$16 \$153 \$8245 VNB sky130_fd_sc_hd__clkbuf_2
X$18692 \$16 \$8353 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18693 \$16 \$8051 \$16 \$153 \$8318 VNB sky130_fd_sc_hd__clkbuf_2
X$18694 \$153 \$8399 \$8318 \$8245 \$8319 \$8288 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$18695 \$153 \$8319 \$8288 \$8287 \$8318 \$8245 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$18696 \$153 \$8318 \$8288 \$8400 \$8319 \$8245 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$18697 \$16 \$8050 \$16 \$153 \$7792 VNB sky130_fd_sc_hd__clkbuf_2
X$18699 \$16 \$7656 \$16 \$153 \$8109 VNB sky130_fd_sc_hd__clkbuf_2
X$18700 \$16 \$7801 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18701 \$16 \$7801 \$16 \$153 \$8111 VNB sky130_fd_sc_hd__clkbuf_2
X$18703 \$16 \$8133 \$16 \$153 \$7880 VNB sky130_fd_sc_hd__clkbuf_2
X$18704 \$16 \$8111 \$8110 \$8109 \$153 \$8134 \$16 VNB sky130_fd_sc_hd__and3b_4
X$18705 \$16 \$7656 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18707 \$16 \$8322 \$16 \$153 \$8220 VNB sky130_fd_sc_hd__clkbuf_2
X$18708 \$16 \$8050 \$16 \$153 \$8354 VNB sky130_fd_sc_hd__clkbuf_2
X$18709 \$16 \$8320 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18712 \$16 \$8051 \$16 \$153 \$8321 VNB sky130_fd_sc_hd__clkbuf_2
X$18713 \$153 \$8401 \$8321 \$8246 \$8225 \$8354 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$18714 \$16 \$8246 \$8354 \$8225 \$8321 \$16 \$153 \$8322 VNB
+ sky130_fd_sc_hd__and4_2
X$18715 \$153 \$8321 \$8354 \$8377 \$8225 \$8246 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$18717 \$153 \$8225 \$8321 \$8323 \$8354 \$8246 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$18718 \$153 \$8225 \$8354 \$8112 \$8321 \$8246 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$18719 \$153 \$7069 \$7375 \$7033 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18720 \$16 \$8391 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18721 \$153 \$8391 \$7131 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$18723 \$153 \$8192 \$7180 \$7033 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18725 \$153 \$153 \$7375 \$8186 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18727 \$16 \$7131 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18728 \$153 \$8018 \$7839 \$8247 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$18729 \$153 \$7116 \$7639 \$7076 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18730 \$153 \$8402 \$8355 \$7131 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18731 \$16 \$8187 \$16 \$153 \$7928 VNB sky130_fd_sc_hd__inv_1
X$18733 \$153 \$8324 \$8018 \$7147 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18734 \$153 \$8324 \$7463 \$7928 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18735 \$153 \$8226 \$8018 \$7174 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18736 \$153 \$8402 \$7208 \$8378 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18737 \$16 \$7147 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18739 \$16 \$7174 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18741 \$153 \$7862 \$9150 \$8248 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$18742 \$153 \$7272 \$7463 \$7076 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18743 \$153 \$8379 \$7180 \$8380 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18745 \$153 \$8135 \$7607 \$8266 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18746 \$16 \$7615 \$16 \$153 \$8199 VNB sky130_fd_sc_hd__clkbuf_2
X$18747 \$153 \$7680 \$7208 \$8266 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18749 \$153 \$8227 \$7862 \$7147 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18750 \$153 \$8381 \$7208 \$8380 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18751 \$16 \$8220 \$16 \$153 \$7939 VNB sky130_fd_sc_hd__inv_1
X$18752 \$153 \$8249 \$7462 \$7939 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18754 \$153 \$8382 \$7462 \$8291 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18756 \$153 \$8325 \$8290 \$7131 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18758 \$153 \$8403 \$8290 \$7133 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18759 \$153 \$8267 \$7375 \$8268 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18761 \$153 \$8191 \$8189 \$7307 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18762 \$16 \$7133 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18763 \$16 \$7307 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18766 \$153 \$8325 \$7208 \$8268 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18767 \$16 \$8044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18769 \$16 \$7353 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18770 \$16 \$7131 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18771 \$153 \$8345 \$8189 \$7353 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18772 \$16 \$8136 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18773 \$16 \$8250 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18774 \$16 \$7464 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18775 \$153 \$8326 \$8189 \$7464 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18776 \$16 \$7307 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18778 \$153 \$8345 \$7375 \$8098 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18779 \$153 \$8326 \$7639 \$8098 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18780 \$16 \$7615 \$16 \$153 \$8032 VNB sky130_fd_sc_hd__clkbuf_2
X$18781 \$153 \$8382 \$8031 \$7377 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18782 \$153 \$7511 \$7639 \$6985 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18783 \$16 \$7377 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18784 \$16 \$6985 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18787 \$16 \$7131 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18788 \$16 \$7464 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18789 \$16 \$6985 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18790 \$153 \$8404 \$8031 \$7464 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18792 \$16 \$7353 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18793 \$153 \$8327 \$8031 \$7353 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18794 \$153 \$8099 \$7463 \$8291 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18795 \$16 \$8291 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18796 \$16 \$8453 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18798 \$16 \$7307 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18801 \$153 \$8252 \$8200 \$7307 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18802 \$16 \$7377 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18803 \$153 \$8346 \$8200 \$7377 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18804 \$153 \$7985 \$7375 \$7882 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18805 \$153 \$8083 \$7208 \$7882 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18808 \$153 \$8328 \$8200 \$7353 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18809 \$16 \$7353 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18810 \$153 \$8084 \$7607 \$7882 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18812 \$16 \$8291 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18813 \$153 \$7863 \$8351 \$8137 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$18814 \$153 \$7916 \$7462 \$7882 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18816 \$153 \$7116 \$7863 \$7464 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18818 \$153 \$8405 \$7863 \$7353 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18819 \$153 \$7960 \$8473 \$8253 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$18820 \$153 \$7369 \$7462 \$7217 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18821 \$16 \$7133 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18822 \$16 \$7147 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18825 \$153 \$8329 \$8330 \$7147 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18826 \$153 \$8383 \$8330 \$7353 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18827 \$16 \$7353 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18828 \$16 \$7131 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18829 \$153 \$7986 \$7462 \$7782 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18830 \$153 \$7680 \$8330 \$7131 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18832 \$16 \$8704 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18833 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$18834 \$16 \$7307 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18835 \$153 \$8269 \$8330 \$7174 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18836 \$153 \$8135 \$8330 \$7307 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18837 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$18838 \$153 \$7584 \$7376 \$7763 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18841 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$18843 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$18844 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$18845 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$18846 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$18847 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$18848 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$18849 \$153 \$2968 \$2643 \$1980 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18851 \$153 \$2109 \$3010 \$1980 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18852 \$153 \$2807 \$1943 \$2785 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18853 \$16 \$1980 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18854 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$18856 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$18857 \$153 \$2845 \$1792 \$2785 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18858 \$16 \$1658 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18859 \$153 \$2969 \$3010 \$1942 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18861 \$16 \$1390 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18862 \$153 \$2736 \$2064 \$2785 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18863 \$153 \$2670 \$3010 \$1795 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18864 \$16 \$1942 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18865 \$16 \$1311 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18867 \$16 \$2932 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18868 \$16 \$1390 \$2932 \$2924 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$18869 \$153 \$2643 \$1311 \$2924 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$18870 \$16 \$1480 \$16 \$153 \$2110 VNB sky130_fd_sc_hd__inv_1
X$18872 \$153 \$3010 \$1595 \$2970 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$18873 \$153 \$2937 \$1815 \$2884 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18875 \$16 \$1795 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18878 \$16 \$2006 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18879 \$153 \$2848 \$2901 \$1795 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18880 \$153 \$2885 \$2901 \$2006 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18881 \$16 \$1795 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18882 \$16 \$1480 \$2932 \$2970 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$18883 \$16 \$981 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18885 \$153 \$2727 \$2901 \$1980 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18886 \$16 \$2932 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18888 \$153 \$2850 \$2901 \$1658 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18889 \$153 \$3011 \$1792 \$2886 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18890 \$16 \$1658 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18891 \$16 \$1980 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18893 \$16 \$1404 \$2932 \$3012 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$18894 \$16 \$2006 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18895 \$153 \$2971 \$2887 \$2006 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18896 \$16 \$2932 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18898 \$153 \$3013 \$2887 \$2180 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18899 \$153 \$2972 \$2887 \$2024 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18900 \$153 \$2971 \$1943 \$3014 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18901 \$153 \$2972 \$2210 \$3014 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18904 \$16 \$2024 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18905 \$16 \$1013 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18907 \$153 \$2853 \$2887 \$1795 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18908 \$16 \$2180 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18909 \$153 \$2938 \$2887 \$1942 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18910 \$153 \$2938 \$2064 \$3014 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18911 \$16 \$1942 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18912 \$16 \$1795 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18914 \$16 \$1291 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18915 \$16 \$1348 \$16 \$153 \$3014 VNB sky130_fd_sc_hd__inv_1
X$18916 \$16 \$1576 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18917 \$16 \$1348 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18918 \$153 \$2939 \$2646 \$2024 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18919 \$16 \$2006 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18920 \$153 \$2854 \$2646 \$1942 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18921 \$16 \$2024 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18922 \$16 \$1795 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18924 \$153 \$2939 \$2210 \$2586 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18925 \$16 \$1594 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18927 \$153 \$2973 \$2646 \$1687 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18928 \$16 \$1942 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18929 \$153 \$2973 \$1792 \$2586 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18930 \$153 \$3038 \$1943 \$3015 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18931 \$153 \$2942 \$2704 \$2180 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18933 \$16 \$1687 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18935 \$153 \$3016 \$1792 \$3015 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18936 \$153 \$2855 \$2704 \$2024 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18937 \$16 \$1264 \$2647 \$3039 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$18938 \$153 \$2990 \$2704 \$1687 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18939 \$16 \$1551 \$2647 \$2941 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$18940 \$16 \$2024 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18943 \$153 \$2940 \$2009 \$3015 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18944 \$153 \$3017 \$1139 \$2941 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$18945 \$153 \$2942 \$2252 \$2671 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18946 \$153 \$2990 \$1792 \$2671 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18947 \$153 \$2974 \$2933 \$2024 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18948 \$16 \$1980 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18951 \$153 \$2943 \$2933 \$1795 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18952 \$16 \$2024 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18953 \$16 \$1942 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18954 \$16 \$1687 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18955 \$153 \$2975 \$2933 \$1687 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18956 \$153 \$2740 \$2009 \$2671 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18957 \$16 \$1795 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18958 \$153 \$2888 \$2933 \$2180 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18961 \$153 \$2976 \$2933 \$2006 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18963 \$153 \$2976 \$1943 \$2889 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18964 \$16 \$2006 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18966 \$16 \$1480 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18967 \$16 \$1658 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18968 \$153 \$2977 \$2933 \$1658 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18970 \$16 \$1390 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18972 \$16 \$1508 \$2647 \$3018 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$18973 \$16 \$1311 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18974 \$153 \$3019 \$2933 \$1980 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18975 \$153 \$2943 \$1815 \$2889 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18976 \$16 \$2195 \$16 \$153 \$2650 VNB sky130_fd_sc_hd__clkbuf_2
X$18977 \$153 \$2977 \$1547 \$2889 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18978 \$16 \$1508 \$16 \$153 \$2634 VNB sky130_fd_sc_hd__inv_1
X$18980 \$153 \$2944 \$2650 \$2538 \$2635 \$2674 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$18981 \$16 \$1480 \$2539 \$2902 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$18982 \$153 \$3020 \$1311 \$2934 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$18983 \$16 \$1390 \$2539 \$2934 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$18985 \$153 \$2978 \$2857 \$1923 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18986 \$16 \$2944 \$16 \$153 \$1496 VNB sky130_fd_sc_hd__clkbuf_2
X$18989 \$153 \$2991 \$3005 \$1923 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18990 \$153 \$2890 \$2857 \$1965 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$18991 \$153 \$3021 \$2184 \$3269 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$18992 \$16 \$2766 \$16 \$153 \$981 VNB sky130_fd_sc_hd__clkbuf_2
X$18993 \$16 \$1480 \$16 \$153 \$2594 VNB sky130_fd_sc_hd__inv_1
X$18994 \$16 \$1390 \$16 \$153 \$3058 VNB sky130_fd_sc_hd__inv_1
X$18997 \$16 \$1965 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$18998 \$153 \$2891 \$2857 \$2089 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19000 \$153 \$2593 \$2857 \$2042 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19001 \$16 \$2089 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19003 \$153 \$3022 \$1471 \$2879 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19004 \$16 \$2042 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19005 \$16 \$1480 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19006 \$153 \$2979 \$2857 \$2043 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19008 \$153 \$2992 \$3020 \$1845 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19009 \$153 \$2498 \$2857 \$1845 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19010 \$16 \$2043 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19011 \$16 \$1845 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19012 \$16 \$2539 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19013 \$16 \$1845 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19014 \$153 \$2893 \$2708 \$1845 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19017 \$153 \$2980 \$2708 \$1805 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19018 \$153 \$2980 \$1703 \$2746 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19019 \$153 \$2981 \$2708 \$2199 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19020 \$16 \$1805 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19021 \$16 \$1845 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19022 \$16 \$1348 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19025 \$153 \$2981 \$2184 \$2746 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19026 \$153 \$2903 \$2708 \$1923 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19027 \$16 \$2199 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19028 \$16 \$1686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19029 \$153 \$2945 \$3006 \$1845 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19030 \$16 \$1923 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19031 \$16 \$1013 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19033 \$16 \$1805 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19035 \$153 \$2903 \$1895 \$2746 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19036 \$16 \$1845 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19037 \$153 \$2993 \$3006 \$2199 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19038 \$153 \$2945 \$1471 \$2925 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19040 \$16 \$2199 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19041 \$153 \$2993 \$2184 \$2925 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19042 \$153 \$2450 \$2359 \$1845 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19044 \$153 \$2946 \$1576 \$3045 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$19045 \$16 \$1923 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19046 \$153 \$2894 \$2946 \$1845 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19048 \$153 \$2994 \$2946 \$2199 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19051 \$153 \$2748 \$2525 \$2043 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19052 \$153 \$2994 \$2184 \$2895 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19053 \$153 \$3023 \$2946 \$2042 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19054 \$16 \$2043 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19055 \$16 \$1845 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19056 \$16 \$3064 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19057 \$153 \$2947 \$1703 \$2895 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19059 \$153 \$3024 \$1171 \$2904 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$19060 \$16 \$3064 \$16 \$153 \$2362 VNB sky130_fd_sc_hd__clkbuf_2
X$19061 \$153 \$2905 \$2597 \$1923 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19063 \$153 \$2948 \$2597 \$2199 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19064 \$16 \$1923 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19065 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$19067 \$153 \$2861 \$1954 \$2346 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19068 \$153 \$3025 \$2184 \$3060 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19069 \$153 \$2948 \$2184 \$2346 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19070 \$16 \$2199 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19072 \$16 \$1508 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19074 \$16 \$1508 \$2347 \$2949 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$19075 \$153 \$3026 \$1703 \$3060 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19076 \$153 \$2950 \$1471 \$3060 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19078 \$153 \$3077 \$1332 \$2949 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$19079 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$19080 \$16 \$2199 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19081 \$153 \$2818 \$1703 \$2637 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19082 \$153 \$2905 \$1895 \$2346 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19083 \$153 \$2880 \$2184 \$2637 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19084 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$19089 \$16 \$1139 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19090 \$153 \$2906 \$1471 \$2637 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19091 \$153 \$2952 \$1139 \$2951 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$19092 \$16 \$1551 \$2347 \$2951 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$19093 \$16 \$1551 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19096 \$153 \$2995 \$1895 \$2926 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19097 \$153 \$2896 \$2952 \$1805 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19099 \$153 \$2995 \$2952 \$1923 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19100 \$16 \$1551 \$16 \$153 \$2926 VNB sky130_fd_sc_hd__inv_1
X$19102 \$153 \$2953 \$2952 \$1845 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19103 \$16 \$2042 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19104 \$16 \$1923 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19105 \$16 \$2043 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19106 \$16 \$2089 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19107 \$153 \$2996 \$2952 \$1965 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19109 \$153 \$2907 \$2952 \$2089 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19110 \$153 \$2996 \$1806 \$2926 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19111 \$153 \$2907 \$2026 \$2926 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19112 \$16 \$3354 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19113 \$16 \$1965 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19114 \$153 \$2750 \$2863 \$2016 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19116 \$16 \$3096 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19118 \$153 \$2953 \$1471 \$2926 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19119 \$16 \$3435 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19121 \$153 \$3098 \$1471 \$2908 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19122 \$153 \$2897 \$2863 \$2105 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19123 \$16 \$2908 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19124 \$16 \$2098 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19125 \$16 \$2016 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19127 \$153 \$2909 \$2863 \$1969 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19128 \$16 \$2908 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19129 \$16 \$2105 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19131 \$153 \$2997 \$2863 \$1756 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19133 \$16 \$2104 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19134 \$153 \$2910 \$2863 \$2104 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19135 \$16 \$1878 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19136 \$16 \$1756 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19137 \$16 \$1879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19141 \$16 \$2166 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19142 \$153 \$3027 \$1868 \$2639 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19143 \$153 \$2910 \$2092 \$2639 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19145 \$16 \$2104 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19146 \$153 \$2821 \$1712 \$2161 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19147 \$153 \$2927 \$2731 \$2104 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19148 \$16 \$1969 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19151 \$16 \$2098 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19152 \$153 \$2927 \$2092 \$2752 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19153 \$153 \$2911 \$1712 \$2752 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19155 \$153 \$2998 \$2731 \$1969 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19156 \$153 \$2912 \$2731 \$2098 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19158 \$153 \$2912 \$1993 \$2752 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19159 \$153 \$2731 \$1760 \$3028 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$19161 \$16 \$2016 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19162 \$153 \$2955 \$2696 \$2016 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19163 \$16 \$2098 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19164 \$16 \$2105 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19165 \$153 \$2999 \$2696 \$1756 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19167 \$16 \$1585 \$2935 \$2954 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$19169 \$153 \$2955 \$1715 \$2627 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19170 \$153 \$2913 \$2092 \$2627 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19171 \$153 \$2999 \$1712 \$2627 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19172 \$16 \$2935 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19174 \$16 \$2104 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19175 \$153 \$2865 \$2796 \$2104 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19176 \$16 \$3198 \$16 \$153 \$2659 VNB sky130_fd_sc_hd__clkbuf_2
X$19178 \$16 \$3198 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19180 \$16 \$1878 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19181 \$16 \$2098 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19183 \$153 \$3062 \$2796 \$2098 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19184 \$153 \$3000 \$2796 \$1878 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19186 \$16 \$901 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19187 \$16 \$2935 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19191 \$16 \$1514 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19192 \$16 \$901 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19194 \$16 \$2105 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19195 \$16 \$1756 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19196 \$153 \$3001 \$2866 \$2105 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19197 \$153 \$2797 \$2866 \$1756 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19198 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$19200 \$16 \$2580 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19201 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$19202 \$16 \$2462 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19203 \$153 \$2866 \$1272 \$2914 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$19205 \$153 \$3029 \$2092 \$2789 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19206 \$153 \$3001 \$2438 \$2789 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19207 \$153 \$2915 \$1558 \$2789 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19208 \$16 \$1272 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19209 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$19210 \$16 \$1878 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19212 \$16 \$1756 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19213 \$16 \$1879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19214 \$153 \$3002 \$2881 \$1756 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19216 \$153 \$2799 \$2881 \$1879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19217 \$153 \$3007 \$2438 \$2790 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19219 \$153 \$2982 \$2881 \$2098 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19220 \$16 \$2098 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19221 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$19223 \$153 \$2982 \$1993 \$2790 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19224 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$19225 \$16 \$815 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19226 \$16 \$2104 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19228 \$16 \$2098 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19229 \$153 \$2801 \$2916 \$2104 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19230 \$153 \$2882 \$2916 \$2098 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19232 \$16 \$1879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19233 \$153 \$3030 \$1613 \$3063 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19234 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$19235 \$16 \$2016 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19236 \$153 \$2928 \$2916 \$2016 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19237 \$16 \$1878 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19238 \$153 \$3003 \$2916 \$1878 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19239 \$153 \$2928 \$1715 \$2791 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19241 \$153 \$3003 \$1868 \$2791 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19243 \$153 \$2956 \$2916 \$2105 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19244 \$16 \$1228 \$2580 \$3051 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$19246 \$153 \$2983 \$2916 \$1756 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19247 \$16 \$2105 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19248 \$16 \$2917 \$16 \$153 \$1566 VNB sky130_fd_sc_hd__clkbuf_2
X$19250 \$153 \$2956 \$2438 \$2791 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19251 \$153 \$2957 \$2916 \$1879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19252 \$153 \$2957 \$1558 \$2791 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19253 \$16 \$1879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19254 \$153 \$3031 \$2271 \$2899 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19255 \$153 \$2958 \$1489 \$2929 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$19257 \$153 \$2870 \$2958 \$2191 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19258 \$16 \$1044 \$1972 \$2929 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$19260 \$153 \$2829 \$2958 \$2031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19262 \$153 \$2959 \$2958 \$2093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19264 \$16 \$2085 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19265 \$153 \$2959 \$2265 \$2899 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19266 \$16 \$2093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19268 \$16 \$1760 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19269 \$16 \$1973 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19270 \$16 \$2031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19271 \$153 \$2961 \$2958 \$2192 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19273 \$16 \$2984 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19274 \$16 \$2960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19275 \$153 \$2962 \$2958 \$1960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19277 \$16 \$2192 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19278 \$16 \$1543 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19279 \$153 \$2962 \$2086 \$2899 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19280 \$153 \$2961 \$2269 \$2899 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19281 \$16 \$2984 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19282 \$153 \$2830 \$2000 \$2613 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19283 \$16 \$2191 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19284 \$153 \$2963 \$2831 \$2191 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19285 \$16 \$1885 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19286 \$16 \$1245 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19289 \$16 \$2031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19290 \$153 \$2963 \$2267 \$2872 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19291 \$16 \$2232 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19292 \$16 \$1933 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19294 \$16 \$1973 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19295 \$153 \$2985 \$2831 \$2031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19296 \$153 \$3008 \$2831 \$1973 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19297 \$153 \$2918 \$2265 \$2872 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19299 \$153 \$2919 \$2086 \$2872 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19300 \$16 \$1860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19301 \$153 \$3008 \$2056 \$2872 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19303 \$153 \$2986 \$2832 \$2192 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19304 \$153 \$2985 \$1936 \$2872 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19305 \$153 \$3032 \$2267 \$2780 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19307 \$16 \$2192 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19308 \$153 \$2987 \$2832 \$2031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19309 \$153 \$2986 \$2269 \$2780 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19310 \$16 \$1272 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19311 \$153 \$2874 \$1272 \$2930 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$19312 \$153 \$3009 \$2271 \$2920 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19315 \$16 \$2462 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19316 \$16 \$2085 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19317 \$16 \$2462 \$2531 \$2930 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$19318 \$153 \$3009 \$2874 \$2085 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19319 \$16 \$2192 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19320 \$153 \$2988 \$2874 \$2192 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19322 \$16 \$2031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19323 \$153 \$2988 \$2269 \$2920 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19326 \$16 \$2085 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19327 \$16 \$1960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19328 \$153 \$2921 \$2874 \$1960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19330 \$153 \$2964 \$2874 \$2031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19331 \$153 \$2921 \$2086 \$2920 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19332 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$19333 \$16 \$815 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19335 \$153 \$2964 \$1936 \$2920 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19337 \$16 \$2984 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19338 \$16 \$2191 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19339 \$153 \$2966 \$2804 \$2191 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19340 \$153 \$2965 \$2056 \$2931 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19341 \$153 \$2922 \$2056 \$2759 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19342 \$16 \$1120 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19343 \$16 \$815 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19346 \$16 \$2093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19347 \$153 \$2966 \$2267 \$2759 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19348 \$153 \$3004 \$2804 \$2093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19349 \$16 \$895 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19350 \$16 \$1303 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19351 \$16 \$1228 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19352 \$153 \$2967 \$2086 \$2759 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19353 \$153 \$3004 \$2265 \$2759 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19354 \$16 \$1228 \$2531 \$2989 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$19355 \$16 \$2085 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19359 \$16 \$2085 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19360 \$16 \$2093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19361 \$153 \$2805 \$2883 \$2085 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19362 \$153 \$2900 \$2883 \$2093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19364 \$16 \$1120 \$16 \$153 \$2642 VNB sky130_fd_sc_hd__inv_1
X$19365 \$153 \$3135 \$2271 \$2923 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19366 \$16 \$2191 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19367 \$16 \$1120 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19371 \$16 \$1228 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19372 \$16 \$1860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19373 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$19374 \$153 \$2806 \$2883 \$1860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19375 \$153 \$3033 \$2267 \$2923 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19376 \$16 \$1973 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19377 \$153 \$3034 \$2000 \$2923 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19378 \$153 \$2877 \$2267 \$2642 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19383 \$16 \$2192 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19384 \$16 \$2031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19385 \$153 \$2618 \$2883 \$2192 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19386 \$153 \$3035 \$2883 \$2031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19388 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$19389 \$153 \$3036 \$2269 \$2923 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19392 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$19393 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$19394 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$19395 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$19396 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$19397 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$19398 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$19400 \$153 \$5437 \$5266 \$5403 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19401 \$153 \$5312 \$5266 \$5245 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19402 \$16 \$5403 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19403 \$153 \$5104 \$5266 \$5736 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19404 \$16 \$5245 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19405 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$19408 \$153 \$5438 \$5266 \$5489 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19409 \$153 \$5312 \$5107 \$5120 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19410 \$153 \$5439 \$5266 \$5404 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19411 \$153 \$5313 \$4706 \$5120 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19413 \$16 \$3692 \$16 \$153 \$5120 VNB sky130_fd_sc_hd__inv_1
X$19415 \$16 \$5181 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19416 \$16 \$5404 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19418 \$16 \$5489 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19419 \$153 \$5344 \$5200 \$5274 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19420 \$153 \$5385 \$5200 \$5404 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19421 \$153 \$5344 \$4706 \$5166 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19422 \$16 \$5404 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19425 \$153 \$5385 \$5177 \$5166 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19426 \$16 \$5274 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19427 \$16 \$5314 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19428 \$153 \$5180 \$5200 \$5736 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19430 \$16 \$3767 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19431 \$153 \$5412 \$5405 \$5166 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19432 \$153 \$5315 \$5107 \$5166 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19433 \$16 \$3841 \$16 \$153 \$5166 VNB sky130_fd_sc_hd__inv_1
X$19436 \$16 \$5736 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19438 \$16 \$5176 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19439 \$16 \$5181 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19440 \$16 \$3778 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19441 \$153 \$5386 \$5240 \$5181 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19442 \$153 \$5275 \$5240 \$5736 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19443 \$16 \$5274 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19444 \$153 \$5227 \$4706 \$5276 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19445 \$16 \$5736 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19447 \$16 \$5176 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19449 \$153 \$5386 \$5174 \$5276 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19450 \$153 \$5372 \$5240 \$5245 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19451 \$16 \$3778 \$16 \$153 \$5276 VNB sky130_fd_sc_hd__inv_1
X$19452 \$153 \$5372 \$5107 \$5276 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19453 \$153 \$5345 \$5107 \$5277 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19454 \$16 \$5245 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19455 \$16 \$4079 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19457 \$153 \$5387 \$5267 \$5736 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19459 \$153 \$5345 \$5267 \$5245 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19460 \$153 \$5413 \$5373 \$5277 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19461 \$16 \$5274 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19462 \$16 \$5181 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19463 \$153 \$5267 \$5183 \$5278 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$19464 \$16 \$5245 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19465 \$16 \$5736 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19468 \$153 \$5414 \$5405 \$5277 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19469 \$16 \$3714 \$16 \$153 \$5277 VNB sky130_fd_sc_hd__inv_1
X$19470 \$16 \$3761 \$5176 \$5346 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$19471 \$153 \$5387 \$5055 \$5277 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19472 \$153 \$5347 \$5095 \$5346 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$19474 \$153 \$5374 \$5347 \$5403 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19476 \$153 \$5182 \$5347 \$5245 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19477 \$153 \$5442 \$5347 \$5518 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19478 \$16 \$5245 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19479 \$16 \$5095 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19481 \$153 \$5279 \$5347 \$5274 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19482 \$16 \$5403 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19483 \$16 \$5518 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19486 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$19487 \$153 \$5415 \$5373 \$5168 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19488 \$16 \$5274 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19490 \$153 \$5375 \$5246 \$5736 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19491 \$153 \$5374 \$5405 \$5168 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19492 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$19493 \$16 \$5736 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19494 \$16 \$5274 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19496 \$153 \$5316 \$5107 \$5337 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19497 \$153 \$5416 \$5405 \$5337 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19498 \$153 \$5361 \$5246 \$5274 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19499 \$153 \$5375 \$5055 \$5337 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19500 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$19501 \$153 \$5280 \$5174 \$5337 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19503 \$16 \$5274 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19505 \$153 \$5417 \$5177 \$5337 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19506 \$153 \$5361 \$4706 \$5337 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19508 \$16 \$4822 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19509 \$153 \$5418 \$4706 \$5517 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19510 \$16 \$5268 \$5152 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$19511 \$16 \$5268 \$5376 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$19512 \$16 \$5268 \$5051 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$19513 \$16 \$3886 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19514 \$16 \$5268 \$4812 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$19515 \$16 \$5269 \$4107 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$19516 \$16 \$5269 \$5388 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$19519 \$16 \$5269 \$4269 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$19520 \$153 \$5461 \$3906 \$5348 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$19521 \$16 \$3907 \$5630 \$5348 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$19522 \$16 \$5269 \$5125 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$19523 \$16 \$5269 \$5349 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$19524 \$16 \$5269 \$5230 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$19525 \$16 \$5106 \$5109 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$19526 \$16 \$5269 \$4179 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$19527 \$16 \$5106 \$5065 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$19528 \$153 \$153 \$5107 \$5203 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19529 \$16 \$5106 \$4943 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$19531 \$16 \$16 \$153 VNB sky130_fd_sc_hd__conb_1
X$19534 \$153 \$153 \$5177 \$5203 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19535 \$16 \$4620 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19536 \$153 \$153 \$5373 \$5203 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19537 \$153 \$153 \$4706 \$5203 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19539 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19540 \$153 \$3710 \$1482 \$5373 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19541 \$153 \$153 \$5055 \$5203 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19544 \$153 \$3839 \$1482 \$5405 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19545 \$16 \$5373 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19546 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19547 \$153 \$3554 \$1482 \$5463 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19548 \$16 \$5405 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19550 \$153 \$5362 \$5406 \$5169 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19551 \$16 \$5477 \$16 \$153 \$3310 VNB sky130_fd_sc_hd__clkbuf_2
X$19554 \$153 \$5317 \$5128 \$5324 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19555 \$153 \$5443 \$5128 \$5338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19556 \$153 \$5317 \$5096 \$5169 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19557 \$16 \$5338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19558 \$16 \$5467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19559 \$153 \$5389 \$5128 \$5478 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19560 \$16 \$5324 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19562 \$153 \$5318 \$5128 \$5566 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19563 \$153 \$5389 \$5390 \$5169 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19564 \$16 \$5232 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19565 \$153 \$5419 \$5287 \$5169 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19566 \$16 \$5566 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19567 \$16 \$5566 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19569 \$153 \$5377 \$5248 \$5338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19570 \$16 \$3660 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19572 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$19573 \$16 \$5469 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19574 \$153 \$5377 \$5209 \$5270 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19575 \$153 \$5249 \$5205 \$5270 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19576 \$16 \$4275 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19577 \$16 \$5232 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19578 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$19579 \$16 \$5338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19580 \$16 \$3692 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19582 \$153 \$5251 \$5096 \$5270 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19585 \$16 \$3841 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19586 \$16 \$5271 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19587 \$153 \$5250 \$5069 \$5270 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19588 \$153 \$5420 \$5390 \$5270 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19590 \$16 \$3841 \$5186 \$5282 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$19591 \$153 \$5421 \$5406 \$5270 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19592 \$153 \$5189 \$5350 \$5232 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19593 \$16 \$5324 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19594 \$16 \$4896 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19597 \$153 \$5206 \$5350 \$5324 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19598 \$16 \$3841 \$16 \$153 \$5013 VNB sky130_fd_sc_hd__inv_1
X$19599 \$16 \$5232 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19600 \$153 \$5363 \$5350 \$5271 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19601 \$153 \$5033 \$5350 \$5338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19603 \$153 \$5363 \$5069 \$5013 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19604 \$16 \$5324 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19605 \$16 \$5338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19607 \$16 \$5271 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19608 \$153 \$5422 \$5406 \$5170 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19609 \$153 \$5190 \$5253 \$5324 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19610 \$153 \$5319 \$5069 \$5170 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19611 \$16 \$5271 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19614 \$153 \$5423 \$5390 \$5170 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19615 \$153 \$5191 \$5253 \$5338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19616 \$16 \$5324 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19617 \$153 \$5231 \$5183 \$5272 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$19618 \$153 \$5320 \$5205 \$5170 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19619 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$19622 \$16 \$5338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19623 \$153 \$5424 \$5287 \$5283 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19624 \$16 \$3714 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19626 \$16 \$5271 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19627 \$153 \$5322 \$5231 \$5271 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19628 \$153 \$5321 \$5205 \$5283 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19629 \$153 \$5207 \$5209 \$5283 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19630 \$153 \$5284 \$5231 \$5324 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19632 \$153 \$5445 \$5231 \$5566 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19634 \$153 \$5208 \$5254 \$5338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19635 \$16 \$5324 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19636 \$16 \$5566 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19637 \$16 \$4107 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19638 \$16 \$3997 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19639 \$153 \$5285 \$5205 \$5171 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19641 \$16 \$5338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19642 \$16 \$3997 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19643 \$153 \$5364 \$5254 \$5324 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19644 \$153 \$5425 \$5390 \$5171 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19645 \$16 \$4246 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19646 \$153 \$5426 \$5519 \$5171 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19647 \$153 \$5364 \$5096 \$5171 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19648 \$16 \$5324 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19651 \$16 \$5271 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19652 \$153 \$5273 \$4246 \$5446 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$19654 \$153 \$5378 \$5273 \$5338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19655 \$153 \$5407 \$3906 \$5447 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$19656 \$16 \$3886 \$16 \$153 \$5286 VNB sky130_fd_sc_hd__inv_1
X$19657 \$16 \$5232 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19658 \$16 \$5338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19662 \$153 \$5391 \$5273 \$5478 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19663 \$153 \$5323 \$5273 \$5324 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19664 \$153 \$5391 \$5390 \$5286 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19665 \$153 \$5323 \$5096 \$5286 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19666 \$16 \$5478 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19667 \$153 \$5392 \$5406 \$5286 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19670 \$16 \$5467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19671 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$19672 \$153 \$5448 \$5407 \$5232 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19673 \$16 \$5324 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19674 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$19675 \$153 \$153 \$5209 \$5155 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19676 \$16 \$5232 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19677 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$19678 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$19679 \$16 \$5519 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19680 \$16 \$5271 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19682 \$153 \$5325 \$5407 \$5324 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19683 \$153 \$5394 \$5407 \$5271 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19684 \$153 \$5325 \$5096 \$5339 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19686 \$153 \$5394 \$5069 \$5339 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19688 \$153 \$3599 \$1482 \$5406 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19689 \$16 \$5406 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19691 \$153 \$5393 \$5209 \$5339 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19692 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19694 \$153 \$5365 \$5110 \$4048 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19695 \$16 \$5625 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19696 \$16 \$3960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19698 \$153 \$5097 \$3788 \$5172 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19700 \$153 \$5211 \$3962 \$5172 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19701 \$153 \$5365 \$3858 \$5172 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19702 \$16 \$4048 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19703 \$153 \$5288 \$3716 \$5172 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19704 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$19705 \$153 \$5110 \$5541 \$5449 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$19707 \$16 \$3814 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19708 \$153 \$4799 \$5452 \$5289 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$19710 \$16 \$4834 \$4881 \$5450 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$19711 \$153 \$5326 \$3651 \$5172 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19712 \$153 \$5212 \$3919 \$5172 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19713 \$16 \$4048 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19714 \$16 \$5351 \$16 \$153 \$5172 VNB sky130_fd_sc_hd__inv_1
X$19715 \$153 \$5352 \$5039 \$4048 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19716 \$153 \$5366 \$5470 \$5340 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19718 \$153 \$5040 \$5039 \$3814 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19719 \$153 \$5290 \$5039 \$3960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19720 \$153 \$5352 \$3858 \$5015 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19721 \$16 \$3960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19722 \$16 \$4196 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19723 \$16 \$5259 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19725 \$16 \$3814 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19726 \$16 \$3889 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19727 \$153 \$5291 \$5041 \$3814 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19729 \$16 \$5259 \$4881 \$5451 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$19730 \$16 \$4048 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19731 \$153 \$5395 \$5041 \$3889 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19733 \$153 \$5367 \$3716 \$5016 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19734 \$153 \$5427 \$3858 \$5016 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19735 \$16 \$5259 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19737 \$16 \$5259 \$16 \$153 \$5016 VNB sky130_fd_sc_hd__inv_1
X$19738 \$16 \$3889 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19739 \$16 \$4139 \$5428 \$5429 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$19740 \$153 \$5327 \$5042 \$3889 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19741 \$16 \$4139 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19742 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$19743 \$153 \$5214 \$3651 \$4951 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19744 \$16 \$5331 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19745 \$16 \$5379 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19746 \$16 \$5331 \$4881 \$5453 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$19747 \$16 \$3960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19748 \$153 \$5192 \$5042 \$3960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19750 \$153 \$5327 \$3962 \$4951 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19751 \$16 \$5017 \$4881 \$5430 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$19752 \$153 \$5292 \$3858 \$4951 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19753 \$153 \$5380 \$4931 \$4048 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19754 \$16 \$3814 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19755 \$16 \$3889 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19757 \$153 \$5293 \$4931 \$3814 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19758 \$153 \$5396 \$4931 \$3960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19759 \$16 \$5017 \$16 \$153 \$4992 VNB sky130_fd_sc_hd__inv_1
X$19760 \$153 \$5380 \$3858 \$4992 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19762 \$153 \$5328 \$4952 \$3889 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19765 \$153 \$5397 \$4952 \$4048 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19766 \$16 \$4048 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19767 \$153 \$5328 \$3962 \$5138 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19768 \$153 \$5397 \$3858 \$5138 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19769 \$153 \$5215 \$3651 \$5138 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19770 \$16 \$4168 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19772 \$16 \$3889 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19773 \$16 \$5353 \$16 \$153 \$5138 VNB sky130_fd_sc_hd__inv_1
X$19774 \$153 \$5455 \$4920 \$3889 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19775 \$153 \$5193 \$4920 \$3814 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19776 \$153 \$5431 \$3858 \$4953 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19777 \$16 \$3814 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19779 \$16 \$3814 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19780 \$16 \$5354 \$16 \$153 \$4953 VNB sky130_fd_sc_hd__inv_1
X$19781 \$16 \$3960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19782 \$153 \$5368 \$5043 \$3814 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19784 \$153 \$5456 \$5043 \$3960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19785 \$153 \$5368 \$3651 \$5139 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19787 \$153 \$5432 \$3858 \$5139 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19789 \$16 \$5400 \$16 \$153 \$5139 VNB sky130_fd_sc_hd__inv_1
X$19790 \$16 \$3889 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19792 \$153 \$5329 \$5112 \$3889 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19794 \$153 \$5408 \$3962 \$5139 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19795 \$153 \$5217 \$3939 \$5113 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19796 \$153 \$5296 \$3716 \$5113 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19797 \$153 \$5433 \$5470 \$5434 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19798 \$153 \$5329 \$3962 \$5113 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19800 \$16 \$5354 \$4724 \$5409 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$19802 \$16 \$5400 \$4724 \$5398 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$19803 \$153 \$5330 \$5112 \$3814 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19804 \$16 \$5482 \$4276 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$19805 \$16 \$5355 \$5381 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$19806 \$16 \$5355 \$4168 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$19807 \$16 \$5435 \$16 \$153 \$5482 VNB sky130_fd_sc_hd__clkbuf_2
X$19808 \$16 \$4048 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19809 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19810 \$16 \$5355 \$4152 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$19811 \$16 \$5355 \$4316 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$19813 \$16 \$1482 \$16 \$153 \$5435 VNB sky130_fd_sc_hd__clkbuf_2
X$19814 \$153 \$5330 \$3651 \$5113 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19815 \$16 \$5435 \$16 \$153 \$5355 VNB sky130_fd_sc_hd__clkbuf_2
X$19816 \$16 \$5483 \$5379 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$19818 \$153 \$5356 \$3986 \$5158 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19819 \$16 \$5140 \$16 \$153 \$5351 VNB sky130_fd_sc_hd__clkbuf_2
X$19820 \$16 \$5297 \$16 \$153 \$5331 VNB sky130_fd_sc_hd__clkbuf_2
X$19821 \$153 \$5236 \$3860 \$4954 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19822 \$153 \$3103 \$1482 \$5074 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19824 \$153 \$3210 \$1482 \$5806 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19825 \$16 \$5355 \$4125 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$19826 \$153 \$4887 \$5480 \$5298 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$19827 \$16 \$5195 \$16 \$153 \$5354 VNB sky130_fd_sc_hd__clkbuf_2
X$19828 \$153 \$5410 \$3893 \$4954 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19829 \$16 \$5045 \$16 \$153 \$4562 VNB sky130_fd_sc_hd__clkbuf_2
X$19832 \$153 \$5332 \$5196 \$3826 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19833 \$153 \$5399 \$5196 \$3898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19834 \$153 \$5399 \$3860 \$5114 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19835 \$153 \$5332 \$3893 \$5114 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19836 \$16 \$4129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19837 \$16 \$3898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19838 \$153 \$5333 \$5196 \$4129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19840 \$153 \$5301 \$5196 \$3691 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19841 \$153 \$5333 \$3986 \$5114 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19842 \$16 \$4129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19843 \$153 \$5302 \$5197 \$4129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19844 \$16 \$5351 \$16 \$153 \$5019 VNB sky130_fd_sc_hd__inv_1
X$19846 \$153 \$5382 \$5197 \$3826 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19848 \$16 \$5579 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19850 \$16 \$3898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19851 \$153 \$5457 \$5197 \$3898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19852 \$153 \$5369 \$5197 \$3691 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19854 \$153 \$5303 \$5543 \$5383 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$19855 \$16 \$5259 \$5116 \$5383 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$19857 \$153 \$5334 \$5303 \$3691 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19859 \$153 \$5341 \$5303 \$4129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19860 \$16 \$3691 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19862 \$16 \$5259 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19863 \$153 \$5341 \$3986 \$5117 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19864 \$16 \$4129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19865 \$16 \$3826 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19866 \$153 \$5357 \$5303 \$3826 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19867 \$153 \$5334 \$3142 \$5117 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19869 \$153 \$5357 \$3893 \$5117 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19871 \$16 \$5400 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19872 \$16 \$3826 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19874 \$153 \$5358 \$5198 \$3826 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19875 \$153 \$5370 \$3860 \$5117 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19876 \$16 \$5331 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19877 \$153 \$5358 \$3893 \$5119 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19878 \$16 \$3898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19879 \$16 \$5400 \$4736 \$5458 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$19880 \$16 \$5331 \$16 \$153 \$5119 VNB sky130_fd_sc_hd__inv_1
X$19881 \$153 \$5305 \$5198 \$3898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19882 \$16 \$3691 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19884 \$153 \$5335 \$5198 \$3691 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19886 \$153 \$5236 \$5163 \$3898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19887 \$153 \$5335 \$3142 \$5119 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19888 \$16 \$3567 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19889 \$153 \$5007 \$3893 \$3567 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19891 \$16 \$3898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19893 \$16 \$3691 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19894 \$16 \$4129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19895 \$153 \$5459 \$5163 \$3691 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19896 \$153 \$5336 \$5163 \$4129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19897 \$16 \$3691 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19898 \$16 \$4016 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19899 \$153 \$4766 \$3565 \$5011 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19900 \$16 \$4129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19902 \$16 \$5353 \$4736 \$5384 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$19903 \$153 \$5356 \$5144 \$4129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19904 \$153 \$5401 \$5144 \$3691 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19905 \$16 \$5353 \$16 \$153 \$5158 VNB sky130_fd_sc_hd__inv_1
X$19907 \$16 \$5354 \$4736 \$5371 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$19908 \$153 \$5238 \$3676 \$5011 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19910 \$153 \$5460 \$5144 \$3826 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19911 \$153 \$5342 \$3860 \$4965 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19912 \$153 \$5199 \$5306 \$5371 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$19913 \$16 \$3826 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19915 \$153 \$5402 \$3986 \$4965 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19917 \$16 \$4129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19918 \$153 \$5402 \$5199 \$4129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19920 \$16 \$5354 \$16 \$153 \$4965 VNB sky130_fd_sc_hd__inv_1
X$19921 \$153 \$5343 \$3893 \$4965 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19922 \$153 \$5359 \$5938 \$5309 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19923 \$16 \$3691 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19925 \$153 \$5436 \$5635 \$5309 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19926 \$153 \$5360 \$5627 \$5309 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19928 \$153 \$5343 \$5199 \$3826 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19929 \$153 \$5342 \$5199 \$3898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19930 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$19931 \$16 \$3898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19933 \$153 \$5411 \$5074 \$5692 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19934 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$19937 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$19938 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$19939 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$19940 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$19941 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$19942 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$19943 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$19944 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$19946 \$153 \$5175 \$5486 \$5181 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19948 \$153 \$5693 \$5710 \$5403 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19949 \$153 \$5662 \$5486 \$5736 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19950 \$16 \$5403 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19953 \$16 \$5736 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19954 \$153 \$5663 \$5486 \$5518 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19956 \$153 \$4705 \$5486 \$5274 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19957 \$153 \$5729 \$5710 \$5274 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19959 \$153 \$5515 \$5463 \$5120 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19960 \$153 \$5710 \$4083 \$5730 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$19961 \$16 \$5274 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19963 \$153 \$5165 \$5486 \$5404 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19964 \$16 \$3638 \$5176 \$5584 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$19965 \$16 \$4162 \$16 \$153 \$5762 VNB sky130_fd_sc_hd__inv_1
X$19967 \$16 \$5176 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19968 \$16 \$5404 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19969 \$16 \$4083 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19970 \$16 \$3660 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19972 \$16 \$4162 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19973 \$16 \$5181 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19975 \$153 \$5664 \$5628 \$5181 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19976 \$153 \$5638 \$5628 \$5404 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19977 \$153 \$5664 \$5174 \$5618 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19978 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$19980 \$153 \$5638 \$5177 \$5618 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19981 \$16 \$5404 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19982 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$19984 \$153 \$5640 \$5628 \$5274 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19985 \$153 \$5639 \$5405 \$5618 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19987 \$153 \$5640 \$4706 \$5618 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19988 \$16 \$4229 \$16 \$153 \$5618 VNB sky130_fd_sc_hd__inv_1
X$19990 \$16 \$4229 \$5712 \$5731 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$19991 \$16 \$4229 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19993 \$16 \$5274 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19994 \$16 \$4229 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19995 \$153 \$5694 \$5641 \$5245 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19996 \$153 \$5642 \$5641 \$5489 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$19997 \$16 \$5489 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$19998 \$153 \$5694 \$5107 \$5619 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$19999 \$16 \$5245 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20001 \$153 \$5642 \$5373 \$5619 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20003 \$16 \$3879 \$5176 \$5561 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$20004 \$16 \$5181 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20005 \$153 \$5733 \$5641 \$5181 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20006 \$16 \$5176 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20007 \$153 \$5643 \$5641 \$5274 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20008 \$16 \$3879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20010 \$16 \$5201 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20011 \$16 \$3879 \$16 \$153 \$5619 VNB sky130_fd_sc_hd__inv_1
X$20013 \$16 \$5720 \$16 \$153 \$5176 VNB sky130_fd_sc_hd__clkbuf_2
X$20014 \$16 \$5274 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20015 \$16 \$5176 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20016 \$153 \$5695 \$5711 \$5245 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20018 \$153 \$5629 \$5711 \$5404 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20019 \$153 \$5695 \$5107 \$5721 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20020 \$16 \$5404 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20023 \$153 \$5629 \$5177 \$5721 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20024 \$16 \$4106 \$5712 \$5562 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$20025 \$153 \$5734 \$5711 \$5403 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20026 \$153 \$5644 \$5711 \$5274 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20027 \$16 \$4106 \$16 \$153 \$5721 VNB sky130_fd_sc_hd__inv_1
X$20028 \$153 \$5442 \$5463 \$5168 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20030 \$153 \$5644 \$4706 \$5721 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20031 \$16 \$3997 \$5712 \$5585 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$20032 \$16 \$5403 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20034 \$16 \$4106 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20035 \$153 \$5586 \$5645 \$5489 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20036 \$16 \$5181 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20037 \$153 \$5620 \$5645 \$5181 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20039 \$16 \$5489 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20040 \$16 \$3997 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20041 \$153 \$5696 \$5645 \$5518 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20042 \$153 \$5620 \$5174 \$5621 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20043 \$16 \$3658 \$16 \$153 \$5621 VNB sky130_fd_sc_hd__inv_1
X$20044 \$153 \$5645 \$3949 \$5646 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$20045 \$153 \$5696 \$5463 \$5621 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20048 \$153 \$5735 \$5461 \$5181 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20049 \$16 \$3658 \$5630 \$5646 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$20050 \$16 \$5181 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20052 \$153 \$5647 \$5405 \$5517 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20053 \$16 \$5403 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20054 \$16 \$3658 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20056 \$16 \$5489 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20057 \$16 \$4494 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20058 \$153 \$5697 \$5461 \$5489 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20060 \$16 \$5245 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20061 \$16 \$3907 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20063 \$153 \$5587 \$5107 \$5517 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20064 \$153 \$5588 \$5463 \$5517 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20065 \$153 \$5697 \$5373 \$5517 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20067 \$153 \$5723 \$5107 \$5722 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20068 \$16 \$5489 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20069 \$153 \$5563 \$5466 \$5245 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20071 \$153 \$5738 \$5466 \$5489 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20072 \$16 \$5245 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20074 \$153 \$5665 \$5466 \$5403 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20075 \$16 \$5181 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20076 \$153 \$5648 \$5466 \$5181 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20078 \$16 \$5403 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20080 \$16 \$4162 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20081 \$153 \$5648 \$5174 \$5464 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20083 \$16 \$4083 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20084 \$16 \$4162 \$5186 \$5698 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$20085 \$16 \$5186 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20086 \$153 \$5548 \$4083 \$5698 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$20087 \$16 \$4162 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20088 \$153 \$5590 \$5406 \$5622 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20089 \$153 \$5666 \$5548 \$5324 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20091 \$153 \$5740 \$5548 \$5338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20092 \$153 \$5443 \$5209 \$5169 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20093 \$153 \$5666 \$5096 \$5622 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20094 \$16 \$4162 \$16 \$153 \$5622 VNB sky130_fd_sc_hd__inv_1
X$20095 \$153 \$5699 \$5548 \$5469 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20098 \$153 \$5667 \$5548 \$5478 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20099 \$153 \$5724 \$5205 \$5622 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20100 \$153 \$5649 \$5520 \$5324 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20101 \$16 \$5469 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20102 \$16 \$3638 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20103 \$16 \$3638 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20105 \$153 \$5667 \$5390 \$5622 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20106 \$16 \$5324 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20108 \$153 \$5668 \$5520 \$5469 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20109 \$153 \$5591 \$5519 \$5622 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20110 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$20111 \$16 \$5469 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20112 \$16 \$4229 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20113 \$153 \$5741 \$5520 \$5478 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20114 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$20116 \$153 \$5565 \$5520 \$5566 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20117 \$16 \$4229 \$5713 \$5742 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$20118 \$16 \$5338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20119 \$16 \$5478 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20120 \$16 \$5566 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20121 \$153 \$5593 \$5406 \$5013 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20122 \$16 \$4178 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20123 \$16 \$4269 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20124 \$153 \$5669 \$4269 \$5650 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$20126 \$16 \$4178 \$5713 \$5650 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$20127 \$153 \$5744 \$5669 \$5271 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20129 \$153 \$5521 \$5390 \$5013 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20130 \$16 \$5467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20132 \$16 \$5271 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20133 \$153 \$5745 \$5669 \$5324 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20134 \$16 \$4479 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20135 \$16 \$5201 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20137 \$153 \$5651 \$5209 \$5623 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20138 \$16 \$3879 \$5186 \$5652 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$20139 \$153 \$5746 \$5669 \$5566 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20140 \$153 \$5653 \$5201 \$5652 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$20141 \$16 \$5324 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20143 \$16 \$5566 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20144 \$153 \$5670 \$5653 \$5338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20145 \$16 \$5186 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20147 \$16 \$3879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20148 \$153 \$5671 \$5653 \$5324 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20149 \$153 \$5522 \$5287 \$5170 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20150 \$16 \$3879 \$16 \$153 \$5595 VNB sky130_fd_sc_hd__inv_1
X$20151 \$16 \$5338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20152 \$16 \$5324 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20155 \$153 \$5672 \$5653 \$5469 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20156 \$153 \$5700 \$5653 \$5271 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20157 \$16 \$5469 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20158 \$153 \$5700 \$5069 \$5595 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20159 \$16 \$5467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20160 \$153 \$5673 \$5125 \$5597 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$20161 \$16 \$5271 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20164 \$16 \$5125 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20165 \$153 \$5747 \$5673 \$5271 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20167 \$16 \$5469 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20168 \$153 \$5598 \$5673 \$5469 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20169 \$153 \$5747 \$5069 \$5726 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20170 \$16 \$5271 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20172 \$153 \$5725 \$5209 \$5726 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20174 \$153 \$5598 \$5287 \$5726 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20176 \$153 \$5748 \$5673 \$5232 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20177 \$153 \$5495 \$5406 \$5171 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20179 \$16 \$5566 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20181 \$153 \$5654 \$5096 \$5726 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20182 \$16 \$5232 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20185 \$153 \$5549 \$3949 \$5674 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$20186 \$16 \$3658 \$5479 \$5674 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$20188 \$153 \$5675 \$5549 \$5232 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20189 \$16 \$3906 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20190 \$153 \$5599 \$5519 \$5286 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20191 \$16 \$3658 \$16 \$153 \$5631 VNB sky130_fd_sc_hd__inv_1
X$20193 \$16 \$5478 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20195 \$16 \$3907 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20196 \$16 \$5232 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20197 \$153 \$5676 \$5549 \$5271 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20198 \$153 \$5567 \$5549 \$5324 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20199 \$153 \$5676 \$5069 \$5631 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20200 \$16 \$5271 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20201 \$16 \$5324 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20202 \$16 \$3658 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20204 \$153 \$5600 \$5407 \$5566 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20207 \$153 \$5878 \$5519 \$5631 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20208 \$153 \$3415 \$1482 \$5500 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20209 \$153 \$5600 \$5519 \$5339 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20210 \$16 \$5566 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20212 \$16 \$5467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20213 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20216 \$153 \$3351 \$1482 \$5795 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20217 \$153 \$5677 \$5407 \$5467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20218 \$153 \$5677 \$5406 \$5339 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20219 \$153 \$5596 \$1482 \$5881 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20221 \$16 \$5714 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20223 \$153 \$5749 \$5632 \$5714 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20224 \$153 \$5678 \$5632 \$5605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20226 \$153 \$153 \$5755 \$5568 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20227 \$16 \$5605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20228 \$16 \$5881 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20229 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$20231 \$153 \$153 \$5775 \$5568 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20232 \$153 \$153 \$5500 \$5568 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20233 \$16 \$3983 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20234 \$16 \$3983 \$16 \$153 \$5568 VNB sky130_fd_sc_hd__clkbuf_2
X$20235 \$16 \$5702 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20236 \$153 \$5701 \$5632 \$5528 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20238 \$153 \$5496 \$5632 \$5702 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20241 \$16 \$4093 \$16 \$153 \$5471 VNB sky130_fd_sc_hd__inv_1
X$20242 \$16 \$5796 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20243 \$16 \$5528 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20245 \$16 \$5528 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20246 \$16 \$5702 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20247 \$153 \$5366 \$5679 \$5702 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20248 \$153 \$5569 \$5679 \$5528 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20249 \$16 \$4093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20250 \$153 \$5701 \$5500 \$5471 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20251 \$16 \$5605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20253 \$16 \$3870 \$16 \$153 \$5340 VNB sky130_fd_sc_hd__inv_1
X$20254 \$153 \$5602 \$5679 \$5605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20255 \$153 \$5751 \$5679 \$5714 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20256 \$153 \$5602 \$5625 \$5340 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20257 \$16 \$3870 \$5428 \$5601 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$20259 \$16 \$5605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20260 \$153 \$5603 \$5655 \$5605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20262 \$153 \$5570 \$5655 \$5714 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20263 \$153 \$5603 \$5625 \$5571 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20264 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$20266 \$16 \$5702 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20267 \$153 \$5497 \$5655 \$5702 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20269 \$16 \$5528 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20271 \$153 \$5572 \$5655 \$5528 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20272 \$16 \$4139 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20273 \$16 \$4126 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20274 \$16 \$3929 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20275 \$16 \$4139 \$16 \$153 \$5571 VNB sky130_fd_sc_hd__inv_1
X$20276 \$16 \$5714 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20277 \$153 \$5680 \$5755 \$5472 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20279 \$153 \$5680 \$5552 \$5714 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20281 \$16 \$5819 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20283 \$16 \$5528 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20284 \$153 \$5703 \$5625 \$5472 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20285 \$153 \$5499 \$5552 \$5528 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20286 \$153 \$5703 \$5552 \$5605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20287 \$16 \$3929 \$16 \$153 \$5472 VNB sky130_fd_sc_hd__inv_1
X$20290 \$16 \$3889 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20291 \$16 \$5605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20292 \$16 \$4047 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20295 \$16 \$5528 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20296 \$16 \$5605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20297 \$153 \$5681 \$5633 \$5605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20298 \$153 \$5553 \$5633 \$5528 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20299 \$16 \$4724 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20301 \$16 \$5353 \$4724 \$5501 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$20303 \$16 \$5473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20306 \$16 \$5702 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20307 \$16 \$5906 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20308 \$153 \$5573 \$5633 \$5702 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20309 \$16 \$5714 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20310 \$153 \$5753 \$5633 \$5714 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20311 \$153 \$5681 \$5625 \$5624 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20312 \$16 \$5605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20313 \$16 \$5856 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20314 \$153 \$5704 \$5656 \$5605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20316 \$153 \$5682 \$5656 \$5702 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20317 \$153 \$5704 \$5625 \$5727 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20319 \$16 \$5528 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20320 \$16 \$4016 \$5906 \$5604 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$20322 \$16 \$5714 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20323 \$153 \$5555 \$5656 \$5528 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20324 \$16 \$4016 \$16 \$153 \$5727 VNB sky130_fd_sc_hd__inv_1
X$20326 \$153 \$5754 \$5656 \$5714 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20327 \$153 \$5657 \$5658 \$5605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20328 \$153 \$5683 \$5658 \$5528 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20330 \$16 \$5605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20332 \$16 \$5702 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20333 \$16 \$5306 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20334 \$153 \$5433 \$5658 \$5702 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20335 \$16 \$3834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20336 \$16 \$5002 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20337 \$16 \$5714 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20338 \$153 \$5705 \$5658 \$5714 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20339 \$153 \$5683 \$5500 \$5434 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20341 \$153 \$5705 \$5755 \$5434 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20342 \$16 \$3834 \$16 \$153 \$5434 VNB sky130_fd_sc_hd__inv_1
X$20344 \$153 \$5684 \$5634 \$5605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20345 \$153 \$5606 \$5634 \$5702 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20346 \$16 \$5482 \$4196 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$20347 \$16 \$5194 \$5306 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$20348 \$16 \$5194 \$4803 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$20350 \$16 \$5194 \$4831 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$20352 \$16 \$4092 \$5906 \$5607 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$20353 \$153 \$5706 \$5634 \$5528 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20354 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20355 \$153 \$3082 \$1482 \$5627 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20356 \$153 \$5706 \$5500 \$5574 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20357 \$153 \$3145 \$1482 \$5635 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20360 \$16 \$3983 \$16 \$153 \$5715 VNB sky130_fd_sc_hd__clkbuf_2
X$20361 \$153 \$153 \$5635 \$5715 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20362 \$153 \$3146 \$1482 \$5938 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20363 \$153 \$153 \$5575 \$5715 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20364 \$153 \$153 \$5938 \$5715 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20366 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20367 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20368 \$16 \$5609 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20370 \$153 \$5685 \$5576 \$5963 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20371 \$16 \$5509 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20372 \$16 \$5575 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20373 \$153 \$5223 \$3565 \$4954 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20374 \$153 \$5685 \$5806 \$5474 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20375 \$16 \$4093 \$16 \$153 \$5474 VNB sky130_fd_sc_hd__inv_1
X$20377 \$16 \$5636 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20378 \$153 \$5608 \$5576 \$5636 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20380 \$153 \$5716 \$5938 \$5474 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20382 \$153 \$5708 \$5635 \$5474 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20383 \$153 \$5608 \$5509 \$5474 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20385 \$153 \$5758 \$5717 \$5636 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20386 \$16 \$5351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20387 \$16 \$5351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20389 \$16 \$4276 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20390 \$16 \$5636 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20391 \$153 \$5610 \$5484 \$5611 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20392 \$153 \$5717 \$4196 \$5531 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$20393 \$153 \$5659 \$5532 \$5636 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20394 \$16 \$3870 \$16 \$153 \$5475 VNB sky130_fd_sc_hd__inv_1
X$20395 \$16 \$4139 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20398 \$16 \$4196 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20399 \$16 \$4047 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20401 \$16 \$3870 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20402 \$16 \$5963 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20403 \$16 \$5223 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20404 \$153 \$5687 \$5532 \$5963 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20405 \$16 \$5718 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20406 \$153 \$5686 \$5532 \$5718 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20407 \$16 \$3929 \$5485 \$5507 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$20408 \$16 \$3929 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20409 \$16 \$5718 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20412 \$153 \$5688 \$5074 \$5614 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20413 \$16 \$5331 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20414 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$20415 \$16 \$5609 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20416 \$153 \$5688 \$5533 \$5609 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20417 \$153 \$5759 \$5533 \$5718 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20418 \$153 \$5613 \$5806 \$5614 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20419 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$20422 \$16 \$5579 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20423 \$153 \$5689 \$5533 \$5579 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20424 \$16 \$5887 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20425 \$153 \$5690 \$5533 \$5887 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20426 \$16 \$4011 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20427 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$20428 \$153 \$5689 \$5484 \$5614 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20430 \$16 \$5799 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20432 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$20433 \$16 \$5636 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20434 \$153 \$5691 \$5578 \$5636 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20435 \$16 \$5963 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20436 \$153 \$5577 \$5578 \$5963 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20437 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$20438 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$20439 \$16 \$5609 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20440 \$153 \$5580 \$5578 \$5609 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20443 \$153 \$5691 \$5509 \$5559 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20444 \$16 \$4152 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20445 \$153 \$5615 \$5484 \$5559 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20446 \$153 \$5637 \$4152 \$5660 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$20448 \$16 \$5786 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20449 \$153 \$5761 \$5637 \$5786 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20451 \$153 \$4836 \$3142 \$3567 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20452 \$16 \$4016 \$5582 \$5660 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$20453 \$153 \$5709 \$5637 \$5887 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20454 \$153 \$5581 \$5637 \$5636 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20457 \$153 \$5709 \$5627 \$5511 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20458 \$153 \$5626 \$5637 \$5609 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20459 \$16 \$4092 \$5582 \$5616 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$20460 \$153 \$5359 \$5560 \$5718 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20461 \$153 \$5626 \$5074 \$5511 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20464 \$16 \$5767 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20466 \$153 \$5661 \$5560 \$5767 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20467 \$16 \$5963 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20468 \$16 \$4092 \$16 \$153 \$5692 VNB sky130_fd_sc_hd__inv_1
X$20469 \$153 \$5513 \$5560 \$5963 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20471 \$153 \$5719 \$5938 \$5692 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20472 \$153 \$5661 \$5575 \$5309 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20474 \$16 \$3834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20476 \$16 \$5786 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20477 \$16 \$5887 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20478 \$153 \$5436 \$5560 \$5786 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20479 \$153 \$5360 \$5560 \$5887 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20480 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$20481 \$153 \$5967 \$5635 \$5692 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20484 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$20485 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$20486 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$20487 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$20488 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$20489 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$20490 \$153 \$8510 \$8331 \$7041 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20491 \$153 \$8639 \$8638 \$8678 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20492 \$153 \$8632 \$8667 \$8580 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20493 \$153 \$8552 \$8331 \$6784 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20496 \$153 \$8680 \$8737 \$8679 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20497 \$153 \$8552 \$6794 \$8384 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20498 \$16 \$8580 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20499 \$153 \$8564 \$8667 \$8724 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20500 \$16 \$7041 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20501 \$16 \$6907 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20502 \$153 \$8532 \$6732 \$8384 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20504 \$153 \$8632 \$8194 \$8678 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20505 \$16 \$6987 \$8577 \$8578 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$20506 \$153 \$8331 \$8167 \$8456 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$20507 \$16 \$8436 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20508 \$16 \$8724 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20509 \$153 \$8722 \$6813 \$8578 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$20510 \$153 \$8511 \$8333 \$7041 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20511 \$16 \$8580 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20513 \$153 \$8174 \$8722 \$8580 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20514 \$153 \$8481 \$6913 \$8206 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20515 \$153 \$8564 \$8457 \$8678 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20516 \$153 \$8207 \$8722 \$8436 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20517 \$16 \$6987 \$16 \$153 \$7816 VNB sky130_fd_sc_hd__inv_1
X$20519 \$153 \$8482 \$6794 \$8206 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20521 \$16 \$7521 \$8577 \$8633 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$20523 \$153 \$8603 \$8533 \$8580 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20524 \$153 \$8693 \$8533 \$8436 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20525 \$153 \$8385 \$6732 \$8036 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20526 \$16 \$8580 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20528 \$153 \$8295 \$6913 \$8036 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20529 \$16 \$6989 \$8577 \$8534 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$20530 \$16 \$8436 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20532 \$153 \$8605 \$8535 \$8436 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20533 \$153 \$8640 \$8535 \$8580 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20535 \$16 \$6989 \$16 \$153 \$8604 VNB sky130_fd_sc_hd__inv_1
X$20536 \$153 \$8640 \$8194 \$8604 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20537 \$153 \$8553 \$8230 \$6784 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20538 \$153 \$8605 \$8209 \$8604 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20540 \$153 \$8681 \$8457 \$8565 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20542 \$153 \$8553 \$6794 \$8208 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20544 \$153 \$8579 \$8668 \$8436 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20545 \$16 \$7041 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20546 \$16 \$6784 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20547 \$153 \$8579 \$8209 \$8565 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20548 \$153 \$8668 \$7335 \$8536 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$20550 \$153 \$8641 \$8668 \$8580 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20552 \$153 \$8606 \$8272 \$6907 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20553 \$153 \$8641 \$8194 \$8565 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20554 \$153 \$8642 \$7399 \$8694 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$20555 \$16 \$6907 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20556 \$153 \$8566 \$8737 \$8513 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20559 \$153 \$8439 \$8272 \$6784 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20560 \$153 \$8643 \$8642 \$8580 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20561 \$153 \$8088 \$6996 \$7772 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20562 \$153 \$8643 \$8194 \$8513 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20563 \$16 \$8580 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20564 \$153 \$8645 \$8669 \$8724 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20567 \$16 \$6935 \$8504 \$8581 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$20568 \$153 \$8669 \$7226 \$8581 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$20570 \$16 \$8436 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20571 \$16 \$6935 \$16 \$153 \$8515 VNB sky130_fd_sc_hd__inv_1
X$20572 \$16 \$8724 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20573 \$153 \$8682 \$8209 \$8515 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20574 \$16 \$7041 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20576 \$16 \$6860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20577 \$153 \$8440 \$8274 \$6784 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20580 \$153 \$8644 \$8194 \$8515 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20581 \$153 \$8645 \$8457 \$8515 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20582 \$153 \$8459 \$6732 \$8196 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20583 \$16 \$6979 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20584 \$153 \$8740 \$7212 \$8695 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$20585 \$16 \$8554 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20586 \$16 \$8121 \$7154 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$20588 \$153 \$8582 \$8209 \$8567 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20589 \$153 \$8670 \$6792 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$20590 \$16 \$8554 \$153 \$8340 \$16 VNB sky130_fd_sc_hd__clkbuf_4
X$20592 \$16 \$8422 \$8503 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$20593 \$16 \$8410 \$7124 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$20594 \$16 \$8410 \$7547 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$20595 \$153 \$8568 \$6907 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$20598 \$153 \$8671 \$6860 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$20599 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20600 \$153 \$8583 \$8610 \$8256 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20601 \$16 \$6915 \$8635 \$8696 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$20602 \$153 \$8634 \$8340 \$6996 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20604 \$153 \$8555 \$8340 \$6732 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20605 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20607 \$153 \$8672 \$8277 \$9097 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20608 \$16 \$8410 \$7659 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$20609 \$153 \$8607 \$8340 \$6749 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20611 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20613 \$153 \$8697 \$8340 \$6913 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20614 \$153 \$8584 \$8614 \$8569 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20615 \$16 \$6749 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20616 \$153 \$8646 \$8744 \$8686 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20618 \$153 \$8570 \$8651 \$8256 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20620 \$16 \$7044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20621 \$153 \$8586 \$6813 \$8585 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$20622 \$153 \$8646 \$8651 \$8569 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20623 \$16 \$6987 \$8635 \$8585 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$20624 \$16 \$8167 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20626 \$16 \$8635 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20627 \$153 \$8683 \$8614 \$8256 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20628 \$153 \$8570 \$8586 \$8686 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20631 \$16 \$6987 \$16 \$153 \$8256 VNB sky130_fd_sc_hd__inv_1
X$20632 \$16 \$8647 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20634 \$153 \$8684 \$8789 \$8256 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20635 \$153 \$8583 \$8586 \$8556 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20636 \$153 \$8954 \$8804 \$8256 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20637 \$16 \$7044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20638 \$16 \$8556 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20639 \$16 \$8686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20641 \$153 \$8648 \$8587 \$8647 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20642 \$153 \$8608 \$8587 \$8556 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20644 \$153 \$8609 \$7659 \$8518 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$20645 \$153 \$8648 \$8614 \$8685 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20646 \$16 \$6989 \$16 \$153 \$8685 VNB sky130_fd_sc_hd__inv_1
X$20648 \$153 \$8608 \$8610 \$8685 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20650 \$153 \$8571 \$8278 \$6916 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20651 \$16 \$7521 \$16 \$153 \$8424 VNB sky130_fd_sc_hd__inv_1
X$20652 \$153 \$8649 \$8609 \$8647 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20653 \$153 \$8571 \$6867 \$8217 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20656 \$16 \$6916 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20657 \$153 \$8649 \$8614 \$8424 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20658 \$153 \$8588 \$8610 \$8424 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20659 \$16 \$8647 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20660 \$153 \$8444 \$8278 \$7044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20661 \$153 \$8650 \$8464 \$8686 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20662 \$153 \$8537 \$6324 \$8217 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20664 \$16 \$7466 \$16 \$153 \$8687 VNB sky130_fd_sc_hd__inv_1
X$20666 \$153 \$8650 \$8651 \$8687 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20667 \$16 \$7044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20669 \$16 \$7399 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20670 \$153 \$8611 \$7399 \$8519 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$20671 \$16 \$7466 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20672 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$20673 \$153 \$8652 \$8610 \$8687 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20676 \$153 \$8653 \$8611 \$8686 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20677 \$153 \$8445 \$8279 \$7060 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20678 \$153 \$8653 \$8651 \$8572 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20679 \$153 \$8589 \$8818 \$8572 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20680 \$16 \$7000 \$16 \$153 \$8572 VNB sky130_fd_sc_hd__inv_1
X$20681 \$16 \$7060 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20683 \$153 \$8612 \$7226 \$8389 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$20685 \$153 \$8654 \$8611 \$8647 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20687 \$153 \$8557 \$7212 \$8414 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$20688 \$153 \$8698 \$8612 \$8686 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20690 \$16 \$7212 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20692 \$16 \$8686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20693 \$16 \$8647 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20694 \$16 \$6935 \$16 \$153 \$8613 VNB sky130_fd_sc_hd__inv_1
X$20696 \$153 \$8655 \$8612 \$8647 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20697 \$153 \$8520 \$8612 \$8556 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20698 \$16 \$8647 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20699 \$153 \$8615 \$8557 \$8686 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20700 \$16 \$6910 \$16 \$153 \$8688 VNB sky130_fd_sc_hd__inv_1
X$20702 \$153 \$8655 \$8614 \$8613 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20703 \$153 \$8615 \$8651 \$8688 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20704 \$153 \$8616 \$8557 \$8556 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20706 \$153 \$8689 \$8557 \$8647 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20708 \$16 \$8556 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20710 \$16 \$8734 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20712 \$153 \$10361 \$6771 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$20713 \$16 \$8647 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20715 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20716 \$153 \$8636 \$8340 \$6324 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20717 \$16 \$10361 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20718 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20720 \$153 \$8689 \$8614 \$8688 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20721 \$153 \$8590 \$8676 \$8126 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20723 \$153 \$8617 \$8340 \$6906 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20724 \$153 \$8674 \$8340 \$6865 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20725 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20729 \$153 \$8558 \$8340 \$7006 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20730 \$153 \$8656 \$8425 \$7387 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20731 \$153 \$8618 \$8425 \$7082 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20732 \$153 \$8656 \$7490 \$8538 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20733 \$16 \$7387 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20735 \$153 \$8591 \$8425 \$7239 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20736 \$16 \$7006 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20737 \$16 \$7239 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20738 \$16 \$7082 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20739 \$153 \$8468 \$7366 \$8538 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20740 \$16 \$8673 \$16 \$153 \$8538 VNB sky130_fd_sc_hd__inv_1
X$20741 \$153 \$8591 \$7482 \$8538 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20742 \$16 \$7387 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20743 \$153 \$8522 \$8426 \$7239 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20745 \$153 \$8559 \$8426 \$7387 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20746 \$153 \$8699 \$8426 \$7082 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20747 \$153 \$8559 \$7490 \$8373 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20748 \$16 \$8619 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20749 \$16 \$8313 \$16 \$153 \$8373 VNB sky130_fd_sc_hd__inv_1
X$20750 \$153 \$8620 \$3454 \$8617 \$8539 \$7995 \$8592 \$8593 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$20752 \$153 \$8620 \$2820 \$8467 \$8619 \$8073 \$8469 \$8593 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$20753 \$16 \$7934 \$16 \$153 \$8593 VNB sky130_fd_sc_hd__clkbuf_2
X$20754 \$16 \$7949 \$16 \$153 \$8620 VNB sky130_fd_sc_hd__clkbuf_2
X$20755 \$16 \$7949 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20757 \$16 \$7934 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20758 \$153 \$8620 \$3772 \$8636 \$8540 \$8675 \$8594 \$8593 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$20760 \$153 \$8620 \$3048 \$8491 \$8524 \$8283 \$8541 \$8593 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$20761 \$153 \$8657 \$8676 \$7994 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20762 \$153 \$8470 \$7482 \$8043 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20764 \$16 \$7239 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20766 \$16 \$7445 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20767 \$153 \$8595 \$8281 \$7129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20768 \$153 \$8427 \$8281 \$7445 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20769 \$16 \$7877 \$16 \$153 \$8280 VNB sky130_fd_sc_hd__clkbuf_2
X$20770 \$16 \$7129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20771 \$16 \$8594 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20772 \$153 \$8768 \$7482 \$8263 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20773 \$16 \$8560 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20776 \$153 \$8542 \$7366 \$8263 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20777 \$16 \$8626 \$16 \$153 \$8263 VNB sky130_fd_sc_hd__inv_1
X$20778 \$153 \$8700 \$8621 \$7029 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20779 \$153 \$8595 \$7215 \$8263 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20780 \$16 \$7328 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20781 \$153 \$8561 \$8621 \$7328 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20782 \$16 \$7029 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20783 \$16 \$7129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20784 \$16 \$8626 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20786 \$16 \$8626 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20787 \$16 \$7445 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20788 \$153 \$8658 \$8621 \$7445 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20789 \$153 \$8561 \$7366 \$8525 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20790 \$153 \$8396 \$6582 \$8222 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20791 \$153 \$8658 \$7327 \$8525 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20792 \$16 \$7067 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20794 \$153 \$8471 \$7066 \$8047 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20795 \$16 \$8624 \$8573 \$8701 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$20796 \$153 \$8659 \$8677 \$7445 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20797 \$16 \$8316 \$8573 \$8526 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$20798 \$16 \$7489 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20800 \$153 \$8596 \$7066 \$8574 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20801 \$16 \$7445 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20802 \$16 \$7129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20803 \$16 \$8428 \$8573 \$8543 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$20804 \$16 \$8702 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20806 \$153 \$8659 \$7327 \$8574 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20807 \$153 \$8597 \$7215 \$8574 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20808 \$16 \$8453 \$8573 \$8703 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$20809 \$153 \$8622 \$8358 \$7129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20811 \$153 \$8598 \$8358 \$7029 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20813 \$16 \$7129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20814 \$16 \$8428 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20815 \$16 \$7029 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20816 \$153 \$8598 \$7066 \$8527 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20817 \$153 \$8622 \$7215 \$8527 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20819 \$16 \$8265 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20820 \$153 \$8690 \$7066 \$8691 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20821 \$16 \$7445 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20822 \$153 \$8623 \$8358 \$7445 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20823 \$16 \$7129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20825 \$16 \$8704 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20828 \$16 \$8705 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20829 \$153 \$8623 \$7327 \$8527 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20830 \$153 \$8497 \$8358 \$7239 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20831 \$153 \$8358 \$8705 \$8625 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$20832 \$16 \$8165 \$8573 \$8625 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$20833 \$153 \$8733 \$8353 \$8706 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$20836 \$16 \$7180 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20837 \$16 \$8545 \$16 \$153 \$8316 VNB sky130_fd_sc_hd__clkbuf_2
X$20838 \$153 \$8528 \$8319 \$8245 \$8318 \$8288 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$20839 \$153 \$8319 \$8318 \$8637 \$8288 \$8245 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$20840 \$16 \$8544 \$16 \$153 \$8624 VNB sky130_fd_sc_hd__clkbuf_2
X$20841 \$16 \$8637 \$16 \$153 \$8428 VNB sky130_fd_sc_hd__clkbuf_2
X$20842 \$16 \$8400 \$16 \$153 \$8359 VNB sky130_fd_sc_hd__clkbuf_2
X$20843 \$153 \$8592 \$8340 \$7180 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20844 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20847 \$153 \$10383 \$7377 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$20848 \$153 \$8469 \$8340 \$7463 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20849 \$16 \$8546 \$16 \$153 \$8673 VNB sky130_fd_sc_hd__clkbuf_2
X$20850 \$16 \$8735 \$8353 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$20851 \$16 \$8735 \$8351 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$20854 \$16 \$8448 \$16 \$153 \$8626 VNB sky130_fd_sc_hd__clkbuf_2
X$20855 \$16 \$8735 \$8285 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$20856 \$16 \$8547 \$16 \$153 \$8313 VNB sky130_fd_sc_hd__clkbuf_2
X$20857 \$16 \$10361 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20858 \$153 \$10361 \$7464 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$20859 \$16 \$8377 \$16 \$153 \$7996 VNB sky130_fd_sc_hd__clkbuf_2
X$20860 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20861 \$153 \$8541 \$8340 \$7376 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20864 \$153 \$8498 \$7463 \$8429 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20865 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20867 \$16 \$7464 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20868 \$153 \$8548 \$8355 \$7377 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20869 \$153 \$8575 \$8355 \$7464 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20870 \$16 \$8673 \$16 \$153 \$8378 VNB sky130_fd_sc_hd__inv_1
X$20871 \$16 \$8673 \$8199 \$8692 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$20874 \$153 \$8575 \$7639 \$8378 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20876 \$153 \$8660 \$8355 \$7353 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20877 \$153 \$8548 \$7462 \$8378 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20879 \$153 \$8660 \$7375 \$8378 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20880 \$16 \$7353 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20881 \$153 \$7956 \$7376 \$7076 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20883 \$153 \$8661 \$8450 \$7353 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20884 \$153 \$8081 \$7180 \$7076 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20885 \$153 \$8599 \$7462 \$8380 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20886 \$16 \$8313 \$16 \$153 \$8380 VNB sky130_fd_sc_hd__inv_1
X$20887 \$16 \$7377 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20888 \$16 \$7667 \$8824 \$8707 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$20890 \$16 \$7464 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20891 \$153 \$8662 \$8450 \$7464 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20892 \$16 \$7131 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20895 \$16 \$7904 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20896 \$16 \$7996 \$8199 \$8600 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$20897 \$153 \$8290 \$8627 \$8600 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$20898 \$153 \$8662 \$7639 \$8380 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20899 \$16 \$7353 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20900 \$16 \$8626 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20901 \$16 \$8626 \$8199 \$8709 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$20903 \$16 \$7464 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20904 \$153 \$8628 \$8290 \$7464 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20906 \$16 \$7307 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20907 \$153 \$8710 \$8290 \$7307 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20908 \$153 \$8403 \$7180 \$8268 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20909 \$153 \$8628 \$7639 \$8268 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20910 \$16 \$7996 \$16 \$153 \$8268 VNB sky130_fd_sc_hd__inv_1
X$20911 \$16 \$7307 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20914 \$153 \$8663 \$8451 \$7307 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20915 \$153 \$8476 \$7376 \$8268 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20917 \$16 \$7131 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20918 \$153 \$8549 \$7376 \$8529 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20919 \$153 \$8663 \$7607 \$8529 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20920 \$153 \$8562 \$8451 \$7131 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20922 \$16 \$7464 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20924 \$153 \$8664 \$8451 \$7464 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20926 \$153 \$8601 \$7375 \$8529 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20927 \$153 \$8664 \$7639 \$8529 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20928 \$153 \$8562 \$7208 \$8529 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20929 \$16 \$7353 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20931 \$16 \$7464 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20932 \$153 \$8563 \$8508 \$7147 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20933 \$153 \$8665 \$8508 \$7464 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20934 \$153 \$8563 \$7463 \$8419 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20935 \$153 \$8665 \$7639 \$8419 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20936 \$16 \$8624 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20937 \$16 \$7307 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20940 \$16 \$7377 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20943 \$153 \$8711 \$8508 \$7307 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20944 \$16 \$7174 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20945 \$153 \$8530 \$8508 \$7174 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20946 \$16 \$8316 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20947 \$16 \$8285 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20948 \$16 \$8453 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20949 \$153 \$8531 \$8285 \$8712 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$20951 \$16 \$8316 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20952 \$16 \$7133 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20954 \$153 \$8550 \$7180 \$8419 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20955 \$153 \$8708 \$8531 \$7307 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20956 \$153 \$9381 \$8531 \$7133 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20957 \$16 \$8316 \$16 \$153 \$8429 VNB sky130_fd_sc_hd__inv_1
X$20958 \$153 \$8327 \$7375 \$8291 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20959 \$16 \$8291 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20961 \$153 \$8100 \$7376 \$8576 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20962 \$153 \$8023 \$7208 \$8291 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20963 \$153 \$8328 \$7375 \$8576 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20964 \$153 \$8420 \$7639 \$8576 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20965 \$153 \$8252 \$7607 \$8576 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20966 \$16 \$8291 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20967 \$16 \$8666 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20968 \$16 \$7498 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20970 \$16 \$8032 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20971 \$16 \$7133 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20972 \$16 \$7147 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20973 \$153 \$8713 \$8602 \$7133 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20974 \$153 \$8629 \$8602 \$7147 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20975 \$153 \$8172 \$7208 \$8576 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20976 \$153 \$8630 \$8602 \$7131 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20978 \$16 \$8428 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20979 \$16 \$7377 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20980 \$153 \$8714 \$8602 \$7377 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20981 \$153 \$8631 \$8602 \$7174 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20983 \$153 \$7683 \$7607 \$7763 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$20984 \$16 \$7174 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20987 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$20988 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$20989 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$20990 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$20991 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$20992 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$20995 \$16 \$7124 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20996 \$16 \$6915 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$20997 \$153 \$8854 \$8667 \$8950 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20998 \$153 \$8639 \$8667 \$8715 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$20999 \$153 \$8736 \$8667 \$9129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21000 \$16 \$8715 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21001 \$16 \$8950 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21002 \$16 \$9129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21005 \$153 \$8826 \$8194 \$8679 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21006 \$153 \$8756 \$8667 \$8436 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21007 \$16 \$9129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21008 \$16 \$6784 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21010 \$153 \$8779 \$8667 \$9026 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21011 \$16 \$6915 \$16 \$153 \$8678 VNB sky130_fd_sc_hd__inv_1
X$21014 \$16 \$6915 \$8577 \$8716 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$21015 \$153 \$8854 \$8912 \$8678 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21016 \$153 \$8667 \$7124 \$8716 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$21017 \$153 \$8799 \$8885 \$8678 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21018 \$16 \$7041 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21019 \$16 \$6988 \$8577 \$8856 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$21020 \$16 \$9129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21021 \$153 \$8725 \$8722 \$9129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21022 \$16 \$8715 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21025 \$153 \$8779 \$8726 \$8678 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21026 \$153 \$8756 \$8209 \$8678 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21027 \$153 \$8757 \$8722 \$8724 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21028 \$153 \$8736 \$8737 \$8678 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21030 \$153 \$8827 \$8737 \$8723 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21032 \$153 \$8693 \$8209 \$8723 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21033 \$153 \$8780 \$8533 \$8715 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21034 \$153 \$8483 \$8533 \$8724 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21035 \$16 \$8715 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21036 \$16 \$8436 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21037 \$153 \$8603 \$8194 \$8723 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21039 \$16 \$8724 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21040 \$153 \$8781 \$8457 \$8604 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21041 \$153 \$8717 \$8726 \$8723 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21042 \$153 \$8782 \$8535 \$8828 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21043 \$16 \$6989 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21045 \$153 \$8738 \$8737 \$8604 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21047 \$153 \$8781 \$8535 \$8724 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21048 \$153 \$8738 \$8535 \$9129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21049 \$16 \$8724 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21050 \$16 \$9129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21051 \$16 \$7973 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21052 \$16 \$6987 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21053 \$153 \$8758 \$8737 \$8565 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21054 \$153 \$8758 \$8668 \$9129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21056 \$153 \$8783 \$8668 \$9026 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21057 \$153 \$8681 \$8668 \$8724 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21058 \$153 \$8783 \$8726 \$8565 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21059 \$16 \$8436 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21060 \$16 \$9026 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21061 \$16 \$9129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21062 \$16 \$8724 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21064 \$16 \$7466 \$16 \$153 \$8565 VNB sky130_fd_sc_hd__inv_1
X$21066 \$16 \$7466 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21067 \$16 \$8580 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21068 \$153 \$8512 \$8642 \$8724 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21069 \$153 \$8566 \$8642 \$9129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21070 \$16 \$8724 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21071 \$16 \$7000 \$8504 \$8694 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$21072 \$16 \$7000 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21073 \$16 \$7399 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21074 \$16 \$8715 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21075 \$16 \$9129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21077 \$153 \$8739 \$8642 \$8436 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21078 \$153 \$8784 \$8642 \$8715 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21079 \$153 \$8739 \$8209 \$8513 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21080 \$153 \$8784 \$8638 \$8513 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21081 \$16 \$7000 \$16 \$153 \$8513 VNB sky130_fd_sc_hd__inv_1
X$21083 \$153 \$8514 \$8669 \$9129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21086 \$153 \$8682 \$8669 \$8436 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21087 \$16 \$9129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21088 \$16 \$8580 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21091 \$153 \$8644 \$8669 \$8580 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21092 \$153 \$8800 \$8726 \$8515 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21094 \$153 \$8829 \$8885 \$8515 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21095 \$153 \$8759 \$8740 \$8580 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21097 \$153 \$8582 \$8740 \$8436 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21098 \$16 \$8580 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21099 \$16 \$6784 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21100 \$16 \$9129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21101 \$153 \$8759 \$8194 \$8567 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21103 \$16 \$6910 \$8504 \$8695 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$21104 \$16 \$6910 \$16 \$153 \$8567 VNB sky130_fd_sc_hd__inv_1
X$21105 \$153 \$8830 \$8885 \$8567 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21106 \$153 \$8741 \$8740 \$9129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21107 \$153 \$8831 \$8726 \$8567 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21108 \$153 \$8741 \$8737 \$8567 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21109 \$16 \$8410 \$8387 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$21111 \$153 \$8832 \$8912 \$8567 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21112 \$153 \$8742 \$8727 \$8256 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21114 \$16 \$6988 \$8635 \$8801 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$21115 \$153 \$8743 \$7124 \$8696 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$21116 \$153 \$8744 \$6888 \$8801 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$21119 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21120 \$153 \$8760 \$8340 \$6794 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21122 \$153 \$8817 \$8744 \$8816 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21124 \$153 \$8584 \$8744 \$8647 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21125 \$16 \$6988 \$16 \$153 \$8569 VNB sky130_fd_sc_hd__inv_1
X$21127 \$16 \$6915 \$16 \$153 \$9097 VNB sky130_fd_sc_hd__inv_1
X$21130 \$16 \$8816 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21132 \$16 \$8898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21133 \$16 \$8647 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21134 \$153 \$8860 \$8744 \$8898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21135 \$16 \$6913 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21136 \$16 \$6996 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21137 \$153 \$8745 \$8744 \$8556 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21138 \$153 \$8785 \$8744 \$8728 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21140 \$153 \$8745 \$8610 \$8569 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21141 \$153 \$8785 \$8818 \$8569 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21142 \$16 \$8686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21143 \$16 \$8556 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21144 \$16 \$6813 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21145 \$16 \$6989 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21146 \$153 \$8683 \$8586 \$8647 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21147 \$153 \$8833 \$8651 \$9097 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21150 \$153 \$8257 \$8586 \$8890 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21151 \$153 \$8366 \$8586 \$8728 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21153 \$153 \$8802 \$8277 \$8424 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21154 \$16 \$6989 \$8635 \$8517 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$21155 \$16 \$8728 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21156 \$153 \$8786 \$8587 \$8728 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21158 \$153 \$8761 \$8587 \$8686 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21159 \$153 \$8761 \$8651 \$8685 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21160 \$16 \$8647 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21161 \$16 \$8686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21162 \$16 \$8556 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21163 \$16 \$6989 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21164 \$16 \$8728 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21165 \$153 \$8746 \$8609 \$8686 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21166 \$16 \$7659 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21169 \$153 \$8786 \$8818 \$8685 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21170 \$16 \$7071 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21171 \$153 \$8465 \$8609 \$8728 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21172 \$16 \$8686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21173 \$16 \$7154 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21174 \$16 \$7521 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21175 \$153 \$8588 \$8609 \$8556 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21177 \$153 \$8746 \$8651 \$8424 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21178 \$153 \$8803 \$8804 \$8424 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21179 \$16 \$8728 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21181 \$153 \$8762 \$8464 \$8728 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21182 \$16 \$8556 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21183 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$21184 \$153 \$8762 \$8818 \$8687 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21186 \$16 \$8686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21187 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$21188 \$16 \$8728 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21190 \$153 \$8763 \$8464 \$8647 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21191 \$153 \$8652 \$8464 \$8556 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21192 \$16 \$8647 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21193 \$153 \$8763 \$8614 \$8687 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21194 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$21197 \$153 \$8589 \$8611 \$8728 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21198 \$153 \$8805 \$8727 \$8687 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21199 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$21200 \$16 \$8686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21201 \$16 \$8728 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21202 \$153 \$8834 \$8727 \$8572 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21204 \$153 \$8747 \$8611 \$8556 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21206 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$21207 \$16 \$8556 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21208 \$153 \$8835 \$8789 \$8572 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21209 \$153 \$8654 \$8614 \$8572 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21210 \$153 \$8748 \$8612 \$8728 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21211 \$153 \$8747 \$8610 \$8572 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21214 \$153 \$8698 \$8651 \$8613 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21215 \$16 \$8728 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21217 \$153 \$8749 \$8612 \$8886 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21218 \$153 \$8748 \$8818 \$8613 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21220 \$153 \$8749 \$8727 \$8613 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21221 \$16 \$8886 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21222 \$16 \$8886 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21223 \$16 \$6910 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21224 \$153 \$8750 \$8277 \$8613 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21226 \$153 \$8790 \$8557 \$8816 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21227 \$153 \$8490 \$6324 \$8260 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21228 \$153 \$8836 \$8727 \$8688 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21230 \$153 \$8616 \$8610 \$8688 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21231 \$16 \$8816 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21232 \$16 \$6867 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21234 \$153 \$8764 \$8557 \$8728 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21235 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21236 \$153 \$8837 \$8789 \$8688 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21237 \$153 \$8806 \$8340 \$7215 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21238 \$16 \$8728 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21239 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21240 \$153 \$8765 \$8340 \$6867 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21242 \$153 \$8764 \$8818 \$8688 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21243 \$153 \$8787 \$8340 \$7327 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21244 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21245 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21246 \$16 \$8838 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21247 \$153 \$8838 \$7445 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$21248 \$16 \$6865 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21249 \$16 \$9869 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21251 \$153 \$9869 \$7129 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$21253 \$153 \$8839 \$7029 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$21254 \$153 \$8729 \$8425 \$7129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21256 \$153 \$8492 \$7327 \$8538 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21258 \$16 \$8673 \$8280 \$8718 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$21259 \$16 \$7344 \$8819 \$8791 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$21260 \$153 \$8425 \$8719 \$8718 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$21261 \$153 \$8861 \$8426 \$7067 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21263 \$153 \$8729 \$7215 \$8538 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21264 \$153 \$8792 \$8426 \$7328 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21265 \$153 \$8494 \$7215 \$8373 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21266 \$16 \$8807 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21267 \$153 \$8792 \$7366 \$8373 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21269 \$153 \$8699 \$7065 \$8373 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21273 \$153 \$8426 \$8820 \$8766 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$21274 \$153 \$8751 \$9252 \$7994 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21275 \$16 \$8313 \$8280 \$8766 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$21276 \$153 \$8620 \$2794 \$8765 \$8821 \$8157 \$8393 \$8593 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$21278 \$153 \$8495 \$7066 \$8043 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21279 \$16 \$8767 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21281 \$153 \$8620 \$3509 \$8674 \$8767 \$7833 \$8730 \$8593 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$21282 \$153 \$8841 \$8676 \$8840 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21283 \$153 \$9148 \$9047 \$7994 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21285 \$153 \$8281 \$8731 \$8720 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$21286 \$16 \$7067 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21288 \$153 \$9099 \$8842 \$7994 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21289 \$153 \$8768 \$8281 \$7239 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21290 \$16 \$8936 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21291 \$153 \$8769 \$8281 \$7067 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21292 \$16 \$9200 \$16 \$153 \$7877 VNB sky130_fd_sc_hd__clkbuf_2
X$21294 \$16 \$7130 \$16 \$153 \$8843 VNB sky130_fd_sc_hd__inv_1
X$21295 \$16 \$8626 \$8280 \$8720 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$21296 \$16 \$8807 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21297 \$16 \$7387 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21298 \$16 \$9200 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21299 \$153 \$8793 \$8621 \$7387 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21300 \$153 \$8752 \$8621 \$7129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21301 \$16 \$7082 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21302 \$153 \$8769 \$6582 \$8263 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21303 \$16 \$7067 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21304 \$16 \$7239 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21306 \$153 \$8795 \$8621 \$7239 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21307 \$153 \$8700 \$7066 \$8525 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21309 \$153 \$8621 \$8702 \$8701 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$21310 \$153 \$8795 \$7482 \$8525 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21311 \$16 \$7877 \$16 \$153 \$8573 VNB sky130_fd_sc_hd__clkbuf_2
X$21313 \$16 \$8624 \$16 \$153 \$8525 VNB sky130_fd_sc_hd__inv_1
X$21314 \$153 \$8796 \$8677 \$7328 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21315 \$153 \$8596 \$8677 \$7029 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21316 \$153 \$8796 \$7366 \$8574 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21317 \$16 \$7239 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21318 \$16 \$7029 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21320 \$153 \$8597 \$8677 \$7129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21321 \$16 \$7328 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21323 \$16 \$7387 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21324 \$16 \$7686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21325 \$16 \$7489 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21327 \$16 \$8453 \$16 \$153 \$8574 VNB sky130_fd_sc_hd__inv_1
X$21328 \$153 \$8809 \$7065 \$8574 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21329 \$153 \$8677 \$8732 \$8703 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$21330 \$16 \$8453 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21331 \$16 \$8453 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21332 \$16 \$8732 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21333 \$16 \$7328 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21334 \$16 \$7029 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21335 \$153 \$8797 \$8733 \$7328 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21337 \$153 \$8690 \$8733 \$7029 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21338 \$153 \$8797 \$7366 \$8691 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21339 \$153 \$8770 \$8733 \$7129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21340 \$16 \$8429 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21341 \$16 \$7387 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21343 \$153 \$8798 \$8733 \$7387 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21345 \$16 \$7445 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21346 \$16 \$8704 \$8573 \$8706 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$21347 \$153 \$8771 \$8733 \$7445 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21348 \$153 \$8798 \$7490 \$8691 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21350 \$153 \$8771 \$7327 \$8691 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21352 \$16 \$8704 \$16 \$153 \$8691 VNB sky130_fd_sc_hd__inv_1
X$21353 \$153 \$8560 \$8340 \$7462 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21354 \$153 \$8594 \$8340 \$7607 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21355 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21357 \$153 \$8734 \$7307 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$21358 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21359 \$16 \$8822 \$7347 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$21362 \$16 \$8822 \$7852 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$21363 \$16 \$8822 \$8794 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$21364 \$16 \$8822 \$8869 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$21365 \$16 \$8822 \$7551 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$21367 \$16 \$8822 \$7668 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$21368 \$16 \$8735 \$8666 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$21370 \$16 \$8735 \$8732 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$21371 \$16 \$8823 \$7686 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$21372 \$16 \$8735 \$8702 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$21373 \$16 \$8823 \$8101 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$21374 \$16 \$8823 \$7915 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$21375 \$16 \$8735 \$8705 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$21377 \$16 \$8823 \$7306 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$21379 \$153 \$8416 \$7353 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$21380 \$16 \$8823 \$8772 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$21381 \$16 \$8823 \$7693 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$21382 \$16 \$8823 \$7614 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$21383 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21384 \$153 \$8393 \$8340 \$7375 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21385 \$153 \$8730 \$8340 \$7639 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21387 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21389 \$16 \$7344 \$8824 \$8870 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$21390 \$153 \$8355 \$8719 \$8692 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$21391 \$153 \$8708 \$7607 \$8429 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21392 \$153 \$8871 \$8904 \$8879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21393 \$16 \$7639 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21394 \$16 \$7208 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21395 \$16 \$7307 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21397 \$16 \$7353 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21398 \$153 \$8753 \$8355 \$7307 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21399 \$16 \$8879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21400 \$16 \$8313 \$8199 \$8810 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$21401 \$153 \$8450 \$8820 \$8810 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$21402 \$153 \$8753 \$7607 \$8378 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21403 \$16 \$7377 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21404 \$153 \$8599 \$8450 \$7377 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21406 \$153 \$8872 \$8922 \$8879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21407 \$153 \$8661 \$7375 \$8380 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21408 \$153 \$8811 \$8996 \$8906 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21409 \$16 \$8879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21410 \$16 \$7307 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21411 \$153 \$8812 \$7668 \$8707 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$21413 \$153 \$8754 \$8450 \$7307 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21414 \$16 \$8313 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21416 \$153 \$8874 \$8794 \$8873 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$21417 \$153 \$8754 \$7607 \$8380 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21418 \$153 \$8963 \$9256 \$8995 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21420 \$153 \$8451 \$8731 \$8709 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$21421 \$16 \$7377 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21422 \$153 \$8773 \$8290 \$7377 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21423 \$16 \$8731 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21424 \$16 \$7996 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21425 \$153 \$8710 \$7607 \$8268 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21426 \$16 \$8627 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21427 \$16 \$7377 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21429 \$153 \$8773 \$7462 \$8268 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21430 \$153 \$8774 \$8451 \$7377 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21431 \$16 \$7667 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21433 \$16 \$8165 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21434 \$16 \$8705 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21435 \$153 \$8774 \$7462 \$8529 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21436 \$16 \$8626 \$16 \$153 \$8529 VNB sky130_fd_sc_hd__inv_1
X$21437 \$16 \$8626 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21438 \$16 \$7353 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21439 \$153 \$8601 \$8451 \$7353 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21440 \$16 \$8032 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21441 \$16 \$7489 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21443 \$16 \$7489 \$8825 \$8875 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$21445 \$16 \$8844 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21446 \$153 \$8478 \$7607 \$8291 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21448 \$16 \$8702 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21449 \$153 \$8508 \$8702 \$8721 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$21450 \$153 \$8845 \$9122 \$8846 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21451 \$153 \$8847 \$8923 \$8846 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21453 \$16 \$8624 \$8032 \$8721 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$21454 \$153 \$8755 \$8508 \$7353 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21455 \$153 \$8848 \$9256 \$8846 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21456 \$16 \$8624 \$16 \$153 \$8419 VNB sky130_fd_sc_hd__inv_1
X$21457 \$153 \$8813 \$7376 \$8291 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21458 \$153 \$8755 \$7375 \$8419 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21460 \$153 \$8814 \$8923 \$8849 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21461 \$153 \$8430 \$8508 \$7377 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21462 \$153 \$8850 \$9256 \$8849 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21463 \$153 \$8711 \$7607 \$8419 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21464 \$16 \$8624 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21465 \$16 \$8032 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21466 \$16 \$7614 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21467 \$153 \$8877 \$7614 \$8876 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$21470 \$16 \$8316 \$8032 \$8712 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$21471 \$16 \$7307 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21473 \$153 \$9798 \$8531 \$7377 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21474 \$153 \$8171 \$7180 \$8576 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21475 \$153 \$8851 \$9122 \$8852 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21476 \$16 \$7377 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21477 \$16 \$7429 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21478 \$16 \$7464 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21480 \$16 \$7353 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21481 \$153 \$8775 \$8531 \$7464 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21482 \$153 \$8878 \$8531 \$7353 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21483 \$153 \$8346 \$7462 \$8576 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21484 \$153 \$8602 \$8666 \$8815 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$21488 \$16 \$7353 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21489 \$153 \$8776 \$8602 \$7353 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21490 \$16 \$8428 \$8032 \$8815 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$21491 \$153 \$8713 \$7180 \$8777 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21492 \$153 \$8629 \$7463 \$8777 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21493 \$16 \$8428 \$16 \$153 \$8777 VNB sky130_fd_sc_hd__inv_1
X$21494 \$16 \$8032 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21495 \$16 \$7464 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21496 \$153 \$8778 \$8602 \$7464 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21499 \$16 \$7498 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21501 \$16 \$8844 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21502 \$16 \$7307 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21503 \$153 \$8881 \$8602 \$7307 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21504 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$21506 \$153 \$7844 \$7462 \$7763 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21507 \$153 \$8853 \$8965 \$8947 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21509 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$21511 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$21512 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$21513 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$21514 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$21515 \$153 \$3284 \$5181 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$21517 \$153 \$6538 \$5405 \$6452 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21518 \$153 \$6602 \$6403 \$5181 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21519 \$16 \$3284 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21520 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$21522 \$16 \$5181 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21523 \$153 \$6602 \$5174 \$6452 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21524 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$21526 \$153 \$6603 \$6403 \$5489 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21527 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$21528 \$153 \$6526 \$6403 \$5404 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21529 \$16 \$5489 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21530 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$21532 \$16 \$4902 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21533 \$16 \$4902 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21534 \$16 \$5404 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21535 \$153 \$6517 \$6397 \$5404 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21536 \$153 \$6661 \$6397 \$5489 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21537 \$16 \$5404 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21538 \$16 \$5489 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21539 \$16 \$5181 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21540 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$21541 \$153 \$6527 \$6397 \$5181 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21544 \$153 \$6662 \$6397 \$5518 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21545 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$21546 \$16 \$5518 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21548 \$153 \$6566 \$5463 \$6260 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21550 \$16 \$5181 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21551 \$153 \$6623 \$6251 \$5181 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21553 \$153 \$6566 \$6251 \$5518 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21555 \$153 \$6623 \$5174 \$6260 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21556 \$16 \$5736 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21557 \$16 \$5518 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21558 \$153 \$6691 \$5373 \$6260 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21559 \$16 \$6784 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21561 \$153 \$6604 \$6406 \$5404 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21563 \$153 \$6663 \$6406 \$5489 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21565 \$153 \$6479 \$6406 \$5518 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21567 \$153 \$6664 \$6406 \$5181 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21569 \$16 \$5518 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21570 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$21571 \$16 \$5181 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21573 \$16 \$5489 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21574 \$153 \$6567 \$6398 \$5736 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21576 \$153 \$6665 \$6398 \$5489 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21577 \$153 \$6499 \$5177 \$6409 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21578 \$16 \$5489 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21580 \$16 \$5181 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21581 \$153 \$6568 \$6398 \$5181 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21582 \$153 \$6567 \$5055 \$6409 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21584 \$153 \$6568 \$5174 \$6409 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21585 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$21586 \$16 \$5518 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21587 \$153 \$6518 \$6280 \$5518 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21588 \$16 \$5181 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21590 \$153 \$6605 \$6280 \$5181 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21591 \$153 \$6605 \$5174 \$6412 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21593 \$153 \$6459 \$6280 \$5404 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21594 \$16 \$5518 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21595 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$21598 \$16 \$3333 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21599 \$16 \$6666 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21600 \$153 \$3333 \$5489 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$21601 \$153 \$6606 \$6280 \$5489 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21602 \$16 \$5404 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21603 \$16 \$5489 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21604 \$153 \$6606 \$5373 \$6412 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21605 \$16 \$5181 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21607 \$153 \$6569 \$6341 \$5181 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21609 \$16 \$6646 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21610 \$153 \$6646 \$3288 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$21611 \$153 \$6569 \$5174 \$6316 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21612 \$153 \$6607 \$6341 \$5518 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21614 \$153 \$6480 \$5405 \$6316 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21616 \$16 \$6647 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21617 \$153 \$6482 \$5055 \$6316 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21618 \$153 \$6647 \$3276 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$21619 \$16 \$5518 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21621 \$16 \$3288 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21623 \$153 \$3288 \$5403 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$21624 \$153 \$6648 \$6732 \$6795 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21625 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$21626 \$16 \$232 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21627 \$153 \$6635 \$7003 \$6695 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21628 \$153 \$6608 \$6399 \$5404 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21631 \$16 \$232 \$16 \$153 \$6667 VNB sky130_fd_sc_hd__clkbuf_2
X$21632 \$153 \$6608 \$5177 \$6177 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21633 \$153 \$6519 \$6399 \$5489 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21635 \$153 \$6528 \$6399 \$5181 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21636 \$16 \$5181 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21639 \$153 \$6609 \$6399 \$5518 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21640 \$16 \$6712 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21641 \$153 \$3096 \$5518 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$21642 \$153 \$6570 \$5406 \$6453 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21643 \$153 \$6571 \$6435 \$5324 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21645 \$16 \$6649 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21647 \$153 \$6649 \$1610 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$21648 \$153 \$6571 \$5096 \$6453 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21650 \$16 \$5324 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21651 \$153 \$6572 \$6435 \$5232 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21652 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$21654 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$21656 \$153 \$6572 \$5205 \$6453 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21657 \$153 \$6668 \$6435 \$5478 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21658 \$153 \$6462 \$5406 \$6414 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21659 \$16 \$5478 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21660 \$16 \$5232 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21661 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$21664 \$153 \$6624 \$6353 \$5566 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21665 \$153 \$6573 \$6353 \$5478 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21666 \$153 \$6624 \$5519 \$6414 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21667 \$153 \$6573 \$5390 \$6414 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21670 \$16 \$6669 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21672 \$153 \$6574 \$6287 \$5232 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21673 \$153 \$6575 \$6287 \$5478 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21674 \$153 \$6574 \$5205 \$6262 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21675 \$153 \$6650 \$6865 \$6695 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21676 \$153 \$6575 \$5390 \$6262 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21677 \$16 \$5232 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21681 \$153 \$6651 \$7003 \$6652 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21683 \$153 \$6464 \$6326 \$5469 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21684 \$153 \$6625 \$6326 \$5232 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21685 \$16 \$5469 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21687 \$16 \$5232 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21690 \$153 \$6576 \$5390 \$6264 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21691 \$16 \$6653 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21692 \$153 \$6653 \$1625 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$21693 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$21694 \$153 \$6529 \$6440 \$5469 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21695 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$21698 \$153 \$6626 \$6440 \$5232 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21699 \$16 \$5324 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21700 \$16 \$5469 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21701 \$153 \$6542 \$5096 \$6357 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21703 \$153 \$6626 \$5205 \$6357 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21704 \$153 \$6543 \$5406 \$6357 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21706 \$16 \$5232 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21709 \$153 \$6577 \$5519 \$6357 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21710 \$16 \$6654 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21711 \$153 \$6654 \$1436 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$21713 \$153 \$6578 \$5390 \$6358 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21714 \$153 \$6530 \$6344 \$5324 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21715 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$21718 \$153 \$6670 \$6344 \$5232 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21720 \$153 \$6579 \$5519 \$6358 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21721 \$16 \$5232 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21722 \$16 \$5324 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21723 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$21724 \$153 \$6483 \$5519 \$6122 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21725 \$153 \$6610 \$6001 \$5232 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21727 \$153 \$6531 \$6001 \$5478 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21728 \$16 \$5232 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21730 \$153 \$6671 \$6034 \$5566 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21731 \$153 \$6610 \$5205 \$6122 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21733 \$153 \$6611 \$6034 \$5467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21735 \$153 \$6672 \$6034 \$5232 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21736 \$16 \$5467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21737 \$153 \$6580 \$5390 \$6291 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21738 \$16 \$5232 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21739 \$16 \$5566 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21740 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$21741 \$153 \$6520 \$6361 \$5478 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21742 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$21744 \$153 \$6612 \$6361 \$5232 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21745 \$153 \$6612 \$5205 \$6416 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21747 \$153 \$6613 \$6361 \$5566 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21748 \$16 \$5232 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21749 \$16 \$5478 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21750 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$21752 \$16 \$3508 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21753 \$153 \$6613 \$5519 \$6416 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21754 \$16 \$5566 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21756 \$153 \$3439 \$5467 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$21757 \$153 \$3200 \$5469 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$21759 \$16 \$3439 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21760 \$16 \$1610 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21761 \$16 \$3243 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21762 \$16 \$3373 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21763 \$16 \$3200 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21764 \$16 \$1775 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21766 \$153 \$6627 \$6642 \$5714 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21767 \$153 \$1610 \$5819 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$21768 \$16 \$5714 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21769 \$16 \$1625 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21771 \$153 \$6614 \$7482 \$5932 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21772 \$153 \$6627 \$5755 \$6556 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21773 \$153 \$6581 \$6582 \$5932 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21775 \$153 \$1625 \$5856 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$21776 \$153 \$6583 \$7066 \$5932 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21779 \$153 \$6467 \$6265 \$5702 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21780 \$153 \$6655 \$5881 \$6556 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21782 \$153 \$6642 \$5541 \$6485 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$21783 \$153 \$6697 \$5500 \$6556 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21784 \$16 \$5351 \$16 \$153 \$6556 VNB sky130_fd_sc_hd__inv_1
X$21785 \$16 \$5714 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21788 \$153 \$6584 \$6332 \$5714 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21789 \$153 \$6636 \$5755 \$6616 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21790 \$16 \$5541 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21791 \$16 \$5819 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21792 \$153 \$6673 \$6698 \$5819 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21793 \$153 \$6584 \$5755 \$6267 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21794 \$16 \$5528 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21796 \$16 \$4834 \$6252 \$6615 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$21797 \$153 \$6757 \$5881 \$6616 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21798 \$16 \$4834 \$16 \$153 \$6616 VNB sky130_fd_sc_hd__inv_1
X$21800 \$153 \$6557 \$6585 \$5528 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21801 \$153 \$6544 \$5470 \$6267 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21802 \$153 \$6586 \$5755 \$6617 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21803 \$153 \$6586 \$6585 \$5714 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21805 \$153 \$6557 \$5500 \$6617 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21806 \$153 \$6545 \$5470 \$6234 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21807 \$153 \$6585 \$4756 \$6510 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$21808 \$153 \$6674 \$6643 \$5819 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21811 \$16 \$4949 \$16 \$153 \$6617 VNB sky130_fd_sc_hd__inv_1
X$21813 \$16 \$5528 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21814 \$16 \$4756 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21815 \$153 \$6675 \$6643 \$5528 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21816 \$153 \$6546 \$5625 \$6234 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21818 \$153 \$6643 \$5379 \$6587 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$21819 \$16 \$5331 \$6252 \$6587 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$21822 \$16 \$5331 \$16 \$153 \$6714 VNB sky130_fd_sc_hd__inv_1
X$21823 \$16 \$5528 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21824 \$16 \$5714 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21825 \$153 \$6644 \$6582 \$6656 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21826 \$16 \$5379 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21828 \$16 \$5819 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21829 \$153 \$6588 \$6511 \$5819 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21830 \$153 \$6628 \$6511 \$5528 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21833 \$153 \$6588 \$6200 \$6558 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21834 \$153 \$6628 \$5500 \$6558 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21835 \$16 \$5017 \$16 \$153 \$6558 VNB sky130_fd_sc_hd__inv_1
X$21836 \$153 \$6512 \$5755 \$6558 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21837 \$16 \$5819 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21838 \$153 \$6532 \$6563 \$5819 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21839 \$16 \$5017 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21840 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$21841 \$16 \$5834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21843 \$153 \$6589 \$6563 \$5834 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21845 \$16 \$5353 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21846 \$153 \$6589 \$5881 \$6533 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21847 \$16 \$5796 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21849 \$16 \$4837 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21850 \$16 \$5714 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21851 \$153 \$6486 \$5625 \$6176 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21852 \$153 \$6559 \$6645 \$5714 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21854 \$16 \$6269 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21855 \$16 \$4837 \$6269 \$6590 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$21856 \$153 \$6559 \$5755 \$6560 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21858 \$16 \$5605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21859 \$153 \$6645 \$4803 \$6590 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$21860 \$153 \$6547 \$5470 \$6176 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21862 \$16 \$4837 \$16 \$153 \$6560 VNB sky130_fd_sc_hd__inv_1
X$21863 \$16 \$5796 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21865 \$153 \$6591 \$6400 \$5796 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21866 \$153 \$6534 \$6400 \$5605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21867 \$153 \$6591 \$5775 \$6455 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21869 \$153 \$6629 \$6400 \$5856 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21870 \$16 \$5400 \$16 \$153 \$6455 VNB sky130_fd_sc_hd__inv_1
X$21872 \$153 \$6592 \$6400 \$5702 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21873 \$153 \$6629 \$5795 \$6455 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21874 \$16 \$5354 \$6269 \$6676 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$21875 \$16 \$5856 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21876 \$153 \$6593 \$5500 \$6535 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21877 \$153 \$6637 \$5625 \$6535 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21878 \$153 \$6618 \$6470 \$5856 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21881 \$16 \$5605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21882 \$153 \$6637 \$6470 \$5605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21884 \$153 \$6488 \$6200 \$6535 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21885 \$153 \$6618 \$5795 \$6535 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21887 \$16 \$5354 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21890 \$16 \$5796 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21891 \$16 \$5528 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21892 \$16 \$5354 \$16 \$153 \$6677 VNB sky130_fd_sc_hd__inv_1
X$21893 \$153 \$6593 \$6470 \$5528 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21894 \$153 \$6678 \$6470 \$5796 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21895 \$153 \$1673 \$5718 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$21896 \$16 \$5480 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21897 \$16 \$4834 \$6216 \$6638 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$21899 \$16 \$5718 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21900 \$153 \$6679 \$5480 \$6638 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$21901 \$153 \$6536 \$6349 \$5718 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21902 \$153 \$6630 \$6679 \$5718 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21905 \$153 \$1544 \$5786 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$21906 \$153 \$6630 \$5938 \$6657 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21907 \$16 \$5351 \$6216 \$6680 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$21908 \$153 \$6491 \$5074 \$6273 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21909 \$153 \$6473 \$6244 \$5609 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21912 \$153 \$6681 \$5541 \$6680 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$21913 \$16 \$5609 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21914 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$21915 \$153 \$6550 \$5635 \$6367 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21917 \$16 \$5963 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21918 \$153 \$6594 \$6244 \$5963 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21919 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$21920 \$16 \$5017 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21923 \$16 \$5017 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21924 \$16 \$5498 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21925 \$153 \$6594 \$5806 \$6367 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21926 \$153 \$6658 \$5484 \$6682 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21927 \$16 \$4949 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21928 \$16 \$5017 \$6216 \$6595 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$21929 \$153 \$6659 \$5938 \$6682 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21930 \$153 \$6619 \$5498 \$6595 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$21931 \$16 \$5017 \$16 \$153 \$6639 VNB sky130_fd_sc_hd__inv_1
X$21933 \$16 \$5579 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21934 \$153 \$6660 \$5938 \$6639 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21935 \$16 \$4756 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21936 \$16 \$4949 \$6216 \$6596 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$21937 \$153 \$6401 \$4756 \$6596 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$21938 \$153 \$6631 \$5379 \$6683 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$21939 \$16 \$5963 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21940 \$153 \$6632 \$6401 \$5963 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21942 \$16 \$5636 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21943 \$153 \$6474 \$5074 \$6047 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21945 \$153 \$6597 \$6401 \$5636 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21947 \$153 \$6632 \$5806 \$6456 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21949 \$16 \$5799 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21950 \$16 \$5331 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21951 \$153 \$6597 \$5509 \$6456 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21953 \$16 \$5331 \$16 \$153 \$6633 VNB sky130_fd_sc_hd__inv_1
X$21954 \$16 \$5609 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21955 \$153 \$6634 \$6401 \$5609 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21956 \$153 \$6391 \$5627 \$6048 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21958 \$153 \$6392 \$5938 \$6456 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21959 \$153 \$6640 \$5799 \$6492 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$21961 \$16 \$5718 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21963 \$16 \$4562 \$6255 \$6598 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$21964 \$153 \$6634 \$5074 \$6456 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21965 \$153 \$6620 \$4609 \$6598 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$21966 \$16 \$5400 \$16 \$153 \$6684 VNB sky130_fd_sc_hd__inv_1
X$21967 \$153 \$6551 \$5074 \$6311 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21968 \$153 \$6393 \$5635 \$6311 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21970 \$153 \$6685 \$6620 \$5887 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21971 \$16 \$4562 \$16 \$153 \$6565 VNB sky130_fd_sc_hd__inv_1
X$21972 \$153 \$6427 \$6308 \$5887 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21973 \$16 \$5887 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21975 \$153 \$6686 \$4803 \$6621 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$21977 \$16 \$4837 \$6255 \$6621 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$21979 \$153 \$6564 \$5938 \$6565 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21980 \$153 \$6687 \$6686 \$5579 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$21981 \$16 \$5579 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21983 \$16 \$4837 \$16 \$153 \$6561 VNB sky130_fd_sc_hd__inv_1
X$21985 \$153 \$6599 \$5938 \$6561 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21986 \$16 \$5354 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21987 \$16 \$5354 \$6255 \$6641 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$21988 \$16 \$4837 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21989 \$16 \$5306 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$21991 \$153 \$6688 \$5306 \$6641 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$21992 \$153 \$5010 \$3986 \$4963 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21993 \$153 \$6562 \$4831 \$6600 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$21995 \$153 \$6622 \$5627 \$6457 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$21997 \$16 \$5354 \$16 \$153 \$6601 VNB sky130_fd_sc_hd__inv_1
X$21998 \$153 \$6689 \$6562 \$5579 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22001 \$153 \$6537 \$6562 \$5963 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22002 \$153 \$6476 \$6562 \$5718 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22003 \$16 \$5963 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22005 \$153 \$6396 \$5575 \$6274 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22007 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$22008 \$16 \$5718 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22009 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$22010 \$16 \$5887 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22011 \$16 \$5786 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22012 \$153 \$6622 \$6562 \$5887 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22013 \$153 \$6690 \$6562 \$5786 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22014 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$22015 \$153 \$6373 \$5635 \$6274 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22018 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$22020 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$22021 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$22022 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$22023 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$22024 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$22025 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$22026 \$153 \$6374 \$6178 \$5736 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22027 \$153 \$6275 \$6178 \$5403 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22030 \$16 \$5403 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22031 \$153 \$6275 \$5405 \$6174 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22032 \$16 \$5736 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22035 \$153 \$6374 \$5055 \$6174 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22037 \$153 \$6352 \$6178 \$5518 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22038 \$153 \$6403 \$5226 \$6375 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$22039 \$16 \$5518 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22040 \$16 \$5226 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22041 \$16 \$4902 \$6051 \$6375 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$22042 \$16 \$6051 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22044 \$16 \$5274 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22046 \$153 \$6338 \$6178 \$5489 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22048 \$153 \$6376 \$6397 \$5274 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22049 \$153 \$6338 \$5373 \$6174 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22050 \$153 \$6376 \$4706 \$6257 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22052 \$153 \$6397 \$5314 \$6339 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$22055 \$16 \$4893 \$6051 \$6339 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$22056 \$16 \$6051 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22057 \$153 \$6404 \$5107 \$6257 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22059 \$153 \$6251 \$5051 \$6276 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$22060 \$16 \$4893 \$16 \$153 \$6257 VNB sky130_fd_sc_hd__inv_1
X$22061 \$16 \$5051 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22062 \$153 \$6340 \$6251 \$5403 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22064 \$153 \$6259 \$6251 \$5245 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22066 \$153 \$6405 \$5177 \$6260 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22067 \$153 \$6277 \$4706 \$6260 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22068 \$16 \$5274 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22069 \$16 \$5245 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22070 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$22071 \$153 \$6340 \$5405 \$6260 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22073 \$153 \$6407 \$6406 \$5274 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22074 \$16 \$5080 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22076 \$153 \$6319 \$5405 \$6315 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22077 \$16 \$5489 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22078 \$153 \$6498 \$5055 \$6315 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22079 \$153 \$6406 \$4939 \$6278 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$22082 \$16 \$4939 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22083 \$153 \$6208 \$5463 \$6043 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22084 \$153 \$6408 \$6398 \$5245 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22085 \$16 \$5404 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22086 \$16 \$6051 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22088 \$16 \$5245 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22089 \$153 \$6398 \$4812 \$6320 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$22090 \$16 \$4621 \$6051 \$6320 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$22091 \$16 \$4621 \$16 \$153 \$6409 VNB sky130_fd_sc_hd__inv_1
X$22094 \$153 \$6377 \$6398 \$5274 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22095 \$153 \$6209 \$5107 \$5993 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22097 \$153 \$6280 \$4973 \$6279 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$22098 \$153 \$6377 \$4706 \$6409 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22101 \$153 \$6410 \$6280 \$5403 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22102 \$153 \$6180 \$5948 \$5489 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22103 \$153 \$6378 \$5055 \$6412 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22104 \$16 \$5489 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22106 \$153 \$6181 \$5948 \$5518 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22107 \$16 \$5403 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22108 \$16 \$4947 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22110 \$16 \$5518 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22111 \$16 \$4947 \$16 \$153 \$6412 VNB sky130_fd_sc_hd__inv_1
X$22112 \$153 \$6411 \$4706 \$6412 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22113 \$16 \$5736 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22114 \$16 \$5026 \$5630 \$6321 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$22115 \$153 \$6341 \$5109 \$6321 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$22116 \$153 \$3491 \$5274 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$22118 \$16 \$5109 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22120 \$16 \$5274 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22121 \$153 \$6281 \$5177 \$5890 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22122 \$153 \$6322 \$6341 \$5274 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22123 \$153 \$6322 \$4706 \$6316 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22124 \$16 \$3491 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22125 \$16 \$5026 \$16 \$153 \$6316 VNB sky130_fd_sc_hd__inv_1
X$22127 \$16 \$5245 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22128 \$16 \$5274 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22130 \$153 \$6282 \$6120 \$5274 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22131 \$153 \$6261 \$6120 \$5245 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22132 \$153 \$6282 \$4706 \$6044 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22133 \$153 \$6432 \$6120 \$5403 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22135 \$16 \$5489 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22137 \$153 \$6224 \$6120 \$5489 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22139 \$16 \$4822 \$5630 \$6379 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$22140 \$153 \$6399 \$4943 \$6379 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$22141 \$16 \$4631 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22142 \$16 \$5489 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22143 \$153 \$6183 \$6060 \$5489 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22144 \$16 \$4943 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22147 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$22148 \$16 \$5403 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22149 \$153 \$6433 \$4706 \$6177 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22150 \$153 \$6283 \$5177 \$6045 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22151 \$153 \$6413 \$6399 \$5403 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22152 \$153 \$6342 \$5107 \$6177 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22155 \$16 \$4621 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22156 \$153 \$6184 \$6399 \$5736 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22157 \$16 \$4812 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22158 \$153 \$6284 \$5174 \$6045 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22159 \$16 \$4621 \$5900 \$6323 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$22160 \$153 \$6353 \$4812 \$6323 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$22161 \$153 \$6413 \$5405 \$6177 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22164 \$153 \$6435 \$5226 \$6434 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$22165 \$16 \$5900 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22166 \$153 \$6343 \$6121 \$5338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22167 \$16 \$4902 \$16 \$153 \$6453 VNB sky130_fd_sc_hd__inv_1
X$22169 \$153 \$6380 \$6353 \$5324 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22170 \$16 \$5271 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22171 \$16 \$5338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22172 \$16 \$4902 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22174 \$153 \$6343 \$5209 \$6149 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22175 \$16 \$4621 \$16 \$153 \$6414 VNB sky130_fd_sc_hd__inv_1
X$22177 \$16 \$5324 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22178 \$153 \$6437 \$6353 \$5469 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22179 \$16 \$4621 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22180 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$22181 \$153 \$6354 \$6121 \$5566 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22182 \$16 \$5469 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22185 \$153 \$6415 \$6353 \$5271 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22186 \$153 \$6286 \$6353 \$5338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22187 \$153 \$6354 \$5519 \$6149 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22188 \$16 \$5338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22189 \$16 \$5566 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22191 \$16 \$5324 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22193 \$16 \$5271 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22194 \$153 \$6188 \$6287 \$5324 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22196 \$153 \$6355 \$6287 \$5566 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22197 \$16 \$5080 \$16 \$153 \$6262 VNB sky130_fd_sc_hd__inv_1
X$22198 \$153 \$6189 \$5209 \$6262 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22199 \$16 \$4896 \$5900 \$6325 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$22200 \$153 \$6326 \$4939 \$6325 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$22203 \$153 \$7213 \$6324 \$6695 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22205 \$16 \$5900 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22206 \$153 \$6263 \$6326 \$5338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22207 \$153 \$6356 \$6326 \$5271 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22208 \$16 \$4896 \$16 \$153 \$6264 VNB sky130_fd_sc_hd__inv_1
X$22210 \$16 \$5271 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22211 \$16 \$4893 \$5900 \$6381 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$22212 \$16 \$5338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22213 \$153 \$6288 \$5846 \$5566 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22214 \$153 \$6440 \$5314 \$6381 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$22215 \$153 \$6288 \$5519 \$6032 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22216 \$16 \$5900 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22217 \$16 \$5314 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22218 \$16 \$4896 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22219 \$16 \$4893 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22221 \$16 \$5566 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22222 \$153 \$6382 \$6440 \$5271 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22223 \$16 \$4973 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22224 \$16 \$4893 \$16 \$153 \$6357 VNB sky130_fd_sc_hd__inv_1
X$22226 \$16 \$4947 \$5900 \$6327 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$22227 \$153 \$6344 \$4973 \$6327 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$22228 \$153 \$6382 \$5069 \$6357 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22229 \$16 \$5271 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22232 \$16 \$6328 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22233 \$153 \$6383 \$6344 \$5271 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22234 \$16 \$6328 \$16 \$153 \$1485 VNB sky130_fd_sc_hd__clkbuf_2
X$22236 \$16 \$5566 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22237 \$153 \$6289 \$5519 \$5980 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22238 \$153 \$6383 \$5069 \$6358 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22239 \$16 \$4947 \$16 \$153 \$6358 VNB sky130_fd_sc_hd__inv_1
X$22241 \$153 \$6290 \$5929 \$5469 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22242 \$16 \$5271 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22244 \$153 \$6329 \$6344 \$5338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22245 \$153 \$6329 \$5209 \$6358 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22246 \$16 \$5478 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22247 \$16 \$5338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22248 \$153 \$6290 \$5287 \$5852 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22249 \$16 \$5469 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22251 \$153 \$6384 \$6001 \$5467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22253 \$153 \$6359 \$6001 \$5271 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22254 \$153 \$6359 \$5069 \$6122 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22255 \$16 \$5271 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22256 \$16 \$5026 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22258 \$16 \$5467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22259 \$16 \$4943 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22260 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$22261 \$153 \$6360 \$6034 \$5271 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22262 \$16 \$4494 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22264 \$153 \$6330 \$6034 \$5338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22266 \$153 \$6361 \$4943 \$6292 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$22267 \$153 \$6360 \$5069 \$6291 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22268 \$153 \$6385 \$6361 \$5324 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22269 \$16 \$5338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22271 \$153 \$6330 \$5209 \$6291 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22273 \$153 \$6345 \$5406 \$6416 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22274 \$153 \$6385 \$5096 \$6416 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22275 \$153 \$6293 \$6085 \$5232 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22276 \$16 \$5324 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22277 \$16 \$5467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22278 \$16 \$5714 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22280 \$153 \$6417 \$6361 \$5338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22282 \$153 \$6293 \$5205 \$6175 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22283 \$153 \$6294 \$5519 \$6175 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22284 \$16 \$5338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22285 \$16 \$5469 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22286 \$153 \$3587 \$5271 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$22287 \$16 \$5232 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22289 \$153 \$6295 \$6085 \$5324 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22290 \$153 \$6331 \$6265 \$5714 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22291 \$153 \$6295 \$5096 \$6175 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22292 \$153 \$6196 \$6195 \$5796 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22294 \$16 \$3587 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22295 \$16 \$3720 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22296 \$16 \$5324 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22297 \$153 \$6443 \$6200 \$6418 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22298 \$153 \$6331 \$5755 \$6418 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22299 \$153 \$6386 \$6265 \$5834 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22300 \$16 \$5796 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22301 \$16 \$5702 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22302 \$16 \$5819 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22304 \$16 \$5856 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22305 \$153 \$6296 \$6265 \$5856 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22306 \$153 \$6386 \$5881 \$6418 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22307 \$153 \$6214 \$5625 \$6136 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22308 \$153 \$6296 \$5795 \$6418 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22310 \$16 \$4760 \$6252 \$6297 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$22311 \$16 \$4760 \$16 \$153 \$6418 VNB sky130_fd_sc_hd__inv_1
X$22314 \$16 \$5819 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22316 \$16 \$5834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22317 \$153 \$6298 \$6332 \$5819 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22318 \$16 \$5856 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22319 \$153 \$6266 \$6332 \$5856 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22320 \$153 \$6298 \$6200 \$6267 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22322 \$153 \$6362 \$5881 \$6267 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22324 \$153 \$6362 \$6332 \$5834 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22325 \$153 \$6332 \$4759 \$6363 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$22326 \$16 \$4930 \$6252 \$6363 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$22328 \$16 \$5856 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22329 \$153 \$6364 \$6333 \$5856 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22330 \$16 \$5834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22331 \$16 \$4759 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22332 \$16 \$4930 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22335 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$22337 \$153 \$6364 \$5795 \$6234 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22338 \$153 \$6268 \$6333 \$5714 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22340 \$16 \$5834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22341 \$153 \$6334 \$6333 \$5834 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22342 \$16 \$5714 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22345 \$153 \$6365 \$6333 \$5819 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22346 \$153 \$6365 \$6200 \$6234 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22347 \$153 \$6334 \$5881 \$6234 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22348 \$153 \$6419 \$5775 \$6234 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22350 \$16 \$5605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22351 \$153 \$6299 \$6253 \$5714 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22353 \$153 \$6387 \$6253 \$5605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22354 \$153 \$6299 \$5755 \$6421 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22355 \$153 \$6387 \$5625 \$6421 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22356 \$16 \$5714 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22358 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$22359 \$16 \$5856 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22362 \$153 \$6420 \$5775 \$6421 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22363 \$153 \$6346 \$6253 \$5856 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22364 \$153 \$6236 \$5881 \$6421 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22365 \$16 \$4562 \$6269 \$6317 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$22366 \$153 \$6346 \$5795 \$6421 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22367 \$153 \$6253 \$4609 \$6317 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$22370 \$16 \$6269 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22371 \$16 \$4562 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22372 \$16 \$4609 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22373 \$16 \$5856 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22374 \$16 \$6124 \$16 \$153 \$6269 VNB sky130_fd_sc_hd__clkbuf_2
X$22375 \$153 \$6270 \$6238 \$5856 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22376 \$153 \$6347 \$6238 \$5834 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22377 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$22378 \$153 \$6347 \$5881 \$6176 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22380 \$153 \$6201 \$6238 \$5714 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22381 \$153 \$6422 \$5775 \$6176 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22382 \$16 \$5714 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22385 \$153 \$6239 \$6200 \$6176 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22386 \$16 \$5605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22387 \$16 \$5528 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22388 \$153 \$6300 \$6012 \$5528 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22391 \$153 \$6423 \$6400 \$5834 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22392 \$153 \$6348 \$6012 \$5605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22394 \$16 \$5400 \$6269 \$6335 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$22395 \$153 \$6424 \$6400 \$5819 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22397 \$153 \$6400 \$5799 \$6335 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$22398 \$153 \$6348 \$5625 \$5892 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22400 \$153 \$6301 \$6271 \$5834 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22401 \$153 \$6425 \$5470 \$6535 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22403 \$16 \$5856 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22404 \$153 \$6301 \$5881 \$6318 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22405 \$153 \$6240 \$6200 \$6318 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22406 \$153 \$6366 \$6271 \$5702 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22407 \$153 \$6241 \$5795 \$6318 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22408 \$153 \$6242 \$5625 \$6318 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22410 \$16 \$5702 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22411 \$16 \$4784 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22412 \$16 \$5906 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22414 \$16 \$5714 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22415 \$16 \$5528 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22416 \$153 \$6388 \$6271 \$5528 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22417 \$16 \$5796 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22418 \$153 \$6302 \$6271 \$5796 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22419 \$16 \$4830 \$16 \$153 \$6535 VNB sky130_fd_sc_hd__inv_1
X$22420 \$153 \$6302 \$5775 \$6318 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22422 \$16 \$4759 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22424 \$153 \$6388 \$5500 \$6318 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22425 \$16 \$5579 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22426 \$153 \$6254 \$6349 \$5579 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22427 \$153 \$6349 \$4759 \$6272 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$22428 \$16 \$5636 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22429 \$16 \$4930 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22430 \$16 \$4930 \$16 \$153 \$6273 VNB sky130_fd_sc_hd__inv_1
X$22432 \$16 \$4760 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22434 \$16 \$4760 \$6216 \$6303 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$22435 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$22436 \$153 \$6389 \$6349 \$5786 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22438 \$153 \$6304 \$6349 \$5636 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22439 \$153 \$6389 \$5635 \$6273 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22440 \$153 \$6304 \$5509 \$6273 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22442 \$153 \$6447 \$6244 \$5767 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22443 \$16 \$4760 \$16 \$153 \$6367 VNB sky130_fd_sc_hd__inv_1
X$22445 \$16 \$5718 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22446 \$153 \$6215 \$5509 \$6018 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22448 \$16 \$5579 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22450 \$153 \$6019 \$5938 \$5475 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22451 \$153 \$6390 \$6244 \$5579 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22453 \$153 \$6368 \$6244 \$5718 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22454 \$153 \$6390 \$5484 \$6367 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22455 \$153 \$6368 \$5938 \$6367 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22456 \$16 \$5259 \$6216 \$6305 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$22458 \$153 \$6350 \$6206 \$5963 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22460 \$16 \$5767 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22462 \$153 \$6336 \$6206 \$5767 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22463 \$153 \$6336 \$5575 \$6047 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22465 \$153 \$6337 \$6206 \$5718 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22466 \$153 \$6350 \$5806 \$6047 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22469 \$153 \$6337 \$5938 \$6047 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22470 \$153 \$6391 \$6169 \$5887 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22471 \$153 \$6306 \$6169 \$5963 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22472 \$16 \$5887 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22474 \$16 \$5767 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22475 \$153 \$6307 \$6169 \$5767 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22479 \$16 \$4882 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22480 \$16 \$5718 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22481 \$153 \$6392 \$6401 \$5718 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22482 \$153 \$6307 \$5575 \$6048 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22483 \$153 \$6426 \$5627 \$6456 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22484 \$16 \$4781 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22486 \$16 \$5963 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22488 \$16 \$6078 \$16 \$153 \$6255 VNB sky130_fd_sc_hd__clkbuf_2
X$22489 \$16 \$5786 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22490 \$153 \$6393 \$6308 \$5786 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22491 \$153 \$6309 \$6308 \$5963 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22492 \$153 \$6309 \$5806 \$6311 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22493 \$16 \$4882 \$16 \$153 \$6311 VNB sky130_fd_sc_hd__inv_1
X$22494 \$16 \$4882 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22496 \$16 \$5636 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22499 \$16 \$5718 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22500 \$153 \$6394 \$6308 \$5636 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22501 \$16 \$5887 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22502 \$16 \$5786 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22503 \$153 \$6310 \$5910 \$5887 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22504 \$153 \$6394 \$5509 \$6311 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22505 \$16 \$5473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22506 \$16 \$5353 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22507 \$153 \$6427 \$5627 \$6311 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22510 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$22511 \$16 \$5786 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22512 \$16 \$5718 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22513 \$153 \$6369 \$6351 \$5786 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22514 \$153 \$6402 \$6351 \$5718 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22515 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$22516 \$16 \$5353 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22519 \$16 \$4567 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22520 \$16 \$5963 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22521 \$16 \$5579 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22522 \$16 \$5767 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22523 \$153 \$6370 \$6351 \$5579 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22524 \$153 \$6395 \$6351 \$5767 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22525 \$16 \$4567 \$5582 \$6313 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$22527 \$16 \$5767 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22528 \$153 \$6428 \$5806 \$6274 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22530 \$16 \$5579 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22532 \$153 \$6371 \$6256 \$5579 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22533 \$153 \$6396 \$6256 \$5767 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22534 \$16 \$4567 \$16 \$153 \$6274 VNB sky130_fd_sc_hd__inv_1
X$22536 \$153 \$6372 \$6256 \$5609 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22537 \$16 \$5963 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22538 \$16 \$5609 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22539 \$16 \$4567 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22542 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$22544 \$16 \$5636 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22545 \$153 \$6373 \$6256 \$5786 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22546 \$153 \$6429 \$6256 \$5636 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22547 \$153 \$6314 \$5074 \$5895 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22548 \$16 \$5786 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22551 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$22553 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$22554 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$22555 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$22556 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$22559 \$153 \$7077 \$6986 \$6981 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22560 \$153 \$7120 \$6986 \$7041 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22562 \$16 \$6783 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22563 \$153 \$7120 \$6996 \$7078 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22564 \$16 \$6981 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22565 \$16 \$7041 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22568 \$153 \$7246 \$6986 \$6784 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22569 \$16 \$7041 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22570 \$153 \$7135 \$6859 \$6907 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22571 \$153 \$7247 \$6986 \$6979 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22572 \$16 \$6907 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22573 \$16 \$6784 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22574 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$22577 \$153 \$7100 \$6719 \$7078 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22578 \$153 \$7279 \$6986 \$6907 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22579 \$16 \$6979 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22581 \$153 \$6986 \$7124 \$7150 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$22582 \$16 \$6915 \$7233 \$7150 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$22583 \$16 \$6907 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22584 \$16 \$6988 \$7233 \$7101 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$22587 \$16 \$6987 \$7233 \$7102 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$22588 \$16 \$6988 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22590 \$153 \$7281 \$7053 \$6981 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22591 \$153 \$7188 \$7053 \$6792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22592 \$153 \$7151 \$7053 \$6860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22593 \$16 \$6792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22594 \$16 \$6979 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22597 \$153 \$7136 \$6794 \$7137 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22598 \$153 \$7139 \$7320 \$6784 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22599 \$153 \$7188 \$6719 \$7137 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22600 \$153 \$7054 \$6995 \$7137 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22601 \$16 \$6860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22602 \$153 \$7151 \$6732 \$7137 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22605 \$153 \$7248 \$7320 \$6979 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22606 \$153 \$6782 \$8387 \$7138 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$22607 \$153 \$6928 \$6913 \$6980 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22608 \$16 \$6989 \$7233 \$7138 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$22609 \$16 \$6979 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22612 \$153 \$7218 \$7234 \$6783 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22613 \$153 \$7139 \$6794 \$7140 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22614 \$16 \$7041 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22615 \$16 \$8387 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22616 \$16 \$6989 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22617 \$153 \$7218 \$6749 \$7141 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22618 \$153 \$7152 \$6719 \$7141 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22619 \$153 \$7104 \$6995 \$6815 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22620 \$16 \$6783 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22621 \$16 \$7041 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22623 \$153 \$7249 \$7234 \$6979 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22624 \$153 \$6931 \$6913 \$6815 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22625 \$153 \$6751 \$7154 \$7153 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$22626 \$16 \$6979 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22628 \$16 \$6909 \$7158 \$7155 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$22629 \$153 \$7157 \$7235 \$6907 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22631 \$153 \$6752 \$7156 \$7155 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$22632 \$16 \$6907 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22633 \$153 \$6908 \$7399 \$7189 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$22634 \$153 \$7157 \$6913 \$7142 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22635 \$16 \$7000 \$7158 \$7189 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$22636 \$16 \$7156 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22638 \$153 \$6883 \$6794 \$6733 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22639 \$153 \$7121 \$6908 \$6981 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22640 \$153 \$6761 \$6749 \$6733 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22641 \$153 \$7121 \$6930 \$6914 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22642 \$16 \$7000 \$16 \$153 \$6914 VNB sky130_fd_sc_hd__inv_1
X$22643 \$153 \$7219 \$7236 \$6907 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22646 \$153 \$7105 \$6995 \$6914 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22647 \$16 \$6907 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22649 \$16 \$6981 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22651 \$153 \$7220 \$6785 \$6979 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22652 \$153 \$7122 \$6785 \$7041 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22653 \$153 \$7122 \$6996 \$6795 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22655 \$153 \$7106 \$6930 \$6795 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22656 \$153 \$7123 \$6786 \$6979 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22657 \$153 \$7220 \$6995 \$6795 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22658 \$16 \$6979 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22660 \$153 \$6786 \$7165 \$7287 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$22661 \$16 \$6981 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22664 \$153 \$7123 \$6995 \$6857 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22665 \$153 \$6861 \$7212 \$7107 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$22666 \$16 \$6979 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22667 \$16 \$6981 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22668 \$153 \$6968 \$6861 \$6981 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22669 \$16 \$7165 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22670 \$16 \$7072 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22671 \$16 \$16 \$153 VNB sky130_fd_sc_hd__conb_1
X$22674 \$16 \$7212 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22675 \$16 \$7124 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22676 \$153 \$153 \$6930 \$7250 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22677 \$153 \$153 \$6995 \$7250 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22678 \$16 \$7237 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22679 \$16 \$7041 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22680 \$16 \$7288 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22681 \$16 \$6910 \$16 \$153 \$6710 VNB sky130_fd_sc_hd__inv_1
X$22682 \$16 \$7545 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22683 \$16 \$6910 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22685 \$153 \$7108 \$6996 \$6710 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22686 \$153 \$6755 \$7124 \$7190 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$22688 \$16 \$6915 \$6990 \$7190 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$22690 \$153 \$7159 \$7073 \$6797 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22691 \$153 \$7191 \$7073 \$6862 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22692 \$16 \$6797 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22693 \$153 \$7159 \$6906 \$6982 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22694 \$16 \$6862 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22695 \$16 \$7545 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22699 \$153 \$7221 \$6756 \$6982 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22700 \$16 \$6862 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22701 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$22702 \$153 \$7192 \$7073 \$7060 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22704 \$153 \$7222 \$7073 \$6771 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22705 \$16 \$7060 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22707 \$153 \$7222 \$6865 \$6982 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22709 \$16 \$6771 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22710 \$16 \$6813 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22711 \$153 \$6787 \$6813 \$7160 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$22712 \$153 \$6905 \$7006 \$6711 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22713 \$16 \$6987 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22714 \$16 \$6987 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22715 \$153 \$7025 \$6867 \$6695 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22716 \$153 \$7079 \$6787 \$6991 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22718 \$153 \$7213 \$6787 \$7060 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22719 \$153 \$7161 \$6865 \$7382 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22720 \$153 \$7162 \$6755 \$7060 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22721 \$16 \$6991 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22722 \$153 \$7162 \$6324 \$6713 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22724 \$153 \$7193 \$6755 \$7044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22725 \$16 \$7060 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22727 \$16 \$8387 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22728 \$153 \$6869 \$8387 \$7194 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$22729 \$16 \$6989 \$6990 \$7194 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$22730 \$16 \$7044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22731 \$153 \$7125 \$6869 \$6916 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22733 \$16 \$7154 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22734 \$16 \$7044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22736 \$153 \$7223 \$6869 \$7044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22737 \$153 \$7193 \$7006 \$6713 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22738 \$16 \$6916 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22739 \$16 \$7044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22740 \$16 \$6991 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22741 \$153 \$6788 \$7154 \$7195 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$22743 \$16 \$7071 \$7163 \$7195 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$22745 \$153 \$7125 \$6867 \$6652 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22746 \$153 \$7224 \$6870 \$6862 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22748 \$16 \$6862 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22749 \$153 \$7126 \$6870 \$6916 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22750 \$16 \$7502 \$16 \$153 \$6918 VNB sky130_fd_sc_hd__inv_1
X$22752 \$16 \$6916 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22754 \$153 \$7126 \$6867 \$6918 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22755 \$153 \$7224 \$7003 \$6918 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22756 \$153 \$7127 \$6788 \$6991 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22758 \$153 \$7081 \$6788 \$7060 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22759 \$16 \$6991 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22762 \$16 \$6909 \$7163 \$7225 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$22764 \$153 \$7127 \$6992 \$6801 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22765 \$153 \$6789 \$7156 \$7225 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$22766 \$16 \$6909 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22768 \$153 \$7008 \$6789 \$7060 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22769 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$22770 \$16 \$6935 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22771 \$16 \$6754 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22772 \$16 \$7226 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22774 \$16 \$6991 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22775 \$16 \$7060 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22776 \$16 \$6935 \$7163 \$7164 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$22777 \$16 \$7044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22778 \$153 \$7227 \$7238 \$7044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22779 \$153 \$6790 \$7226 \$7164 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$22780 \$16 \$6797 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22782 \$16 \$7072 \$7163 \$7144 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$22784 \$153 \$7252 \$7212 \$7251 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$22787 \$153 \$6791 \$7165 \$7144 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$22788 \$153 \$7227 \$7006 \$7316 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22789 \$16 \$6935 \$16 \$153 \$6805 VNB sky130_fd_sc_hd__inv_1
X$22790 \$16 \$7165 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22792 \$16 \$6916 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22793 \$153 \$7253 \$7327 \$5932 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22794 \$153 \$7196 \$7252 \$6916 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22797 \$16 \$6910 \$16 \$153 \$7254 VNB sky130_fd_sc_hd__inv_1
X$22798 \$153 \$7196 \$6867 \$7254 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22799 \$153 \$7109 \$6992 \$6805 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22800 \$153 \$7228 \$7252 \$6754 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22801 \$153 \$7026 \$6324 \$6805 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22804 \$153 \$7166 \$6324 \$7254 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22805 \$153 \$7228 \$6756 \$7254 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22806 \$153 \$7197 \$7252 \$6797 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22807 \$153 \$7255 \$7252 \$6991 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22808 \$153 \$7214 \$7252 \$6862 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22809 \$16 \$6991 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22811 \$153 \$7197 \$6906 \$7254 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22812 \$16 \$7044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22813 \$16 \$7044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22814 \$153 \$7045 \$7003 \$6919 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22815 \$153 \$6614 \$7013 \$7239 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22816 \$16 \$6862 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22817 \$16 \$7067 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22818 \$16 \$7239 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22820 \$153 \$7010 \$7013 \$7082 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22821 \$153 \$7256 \$7065 \$7296 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22822 \$153 \$7229 \$7215 \$7257 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22824 \$16 \$7239 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22825 \$153 \$7198 \$7014 \$7239 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22826 \$153 \$7046 \$7066 \$7257 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22828 \$153 \$7229 \$7014 \$7129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22829 \$16 \$7129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22831 \$16 \$7082 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22832 \$153 \$7199 \$7014 \$7082 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22833 \$153 \$7198 \$7482 \$7257 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22834 \$153 \$7258 \$7490 \$7257 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22836 \$153 \$7110 \$6582 \$7257 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22838 \$16 \$7328 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22840 \$153 \$7145 \$7065 \$7146 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22841 \$153 \$7028 \$7215 \$7146 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22842 \$153 \$7128 \$6972 \$7029 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22843 \$153 \$7259 \$7490 \$7146 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22846 \$16 \$7239 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22847 \$153 \$7260 \$6972 \$7239 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22848 \$153 \$7128 \$7066 \$7146 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22850 \$153 \$7167 \$6582 \$7146 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22851 \$16 \$7029 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22852 \$16 \$7239 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22853 \$153 \$7261 \$7074 \$7239 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22855 \$16 \$7129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22857 \$153 \$7083 \$7074 \$7129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22859 \$153 \$7084 \$7074 \$7029 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22861 \$153 \$7200 \$7074 \$7067 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22864 \$153 \$7200 \$6582 \$7085 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22865 \$16 \$7067 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22867 \$16 \$7130 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22868 \$16 \$7082 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22869 \$16 \$7129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22870 \$153 \$7088 \$7086 \$7082 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22871 \$16 \$7239 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22872 \$153 \$7168 \$7086 \$7239 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22875 \$153 \$7168 \$7482 \$7112 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22876 \$153 \$7230 \$7086 \$7129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22877 \$153 \$7111 \$6582 \$7112 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22878 \$153 \$7230 \$7215 \$7112 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22879 \$153 \$7201 \$7169 \$7067 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22882 \$153 \$7015 \$7169 \$7029 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22883 \$16 \$7029 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22885 \$16 \$7129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22886 \$153 \$7202 \$7170 \$7129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22887 \$16 \$7239 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22888 \$153 \$7300 \$7170 \$7239 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22890 \$153 \$7203 \$7170 \$7029 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22891 \$153 \$7201 \$6582 \$7317 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22892 \$16 \$7082 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22893 \$153 \$7068 \$7170 \$7082 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22895 \$153 \$7262 \$7215 \$7264 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22898 \$16 \$7129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22900 \$153 \$7263 \$7482 \$7264 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22901 \$153 \$7204 \$7171 \$7067 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22902 \$153 \$7447 \$7327 \$7264 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22903 \$16 \$7067 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22904 \$153 \$7204 \$6582 \$7264 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22905 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$22908 \$16 \$7029 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22909 \$16 \$7328 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22910 \$16 \$7082 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22911 \$153 \$7266 \$7090 \$7328 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22912 \$16 \$7029 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22913 \$153 \$7205 \$7090 \$7082 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22914 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$22915 \$153 \$7113 \$7066 \$7172 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22917 \$16 \$7387 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22921 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$22922 \$16 \$7067 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22923 \$153 \$7304 \$7265 \$7067 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22925 \$153 \$7114 \$6582 \$7172 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22926 \$153 \$7030 \$5470 \$6715 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22927 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$22928 \$16 \$7239 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22929 \$153 \$7305 \$7265 \$7239 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22931 \$153 \$7216 \$7090 \$7239 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22932 \$153 \$6592 \$5470 \$6455 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22933 \$16 \$7239 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22934 \$153 \$6952 \$5625 \$6715 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22935 \$16 \$7267 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22936 \$16 \$7306 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22938 \$153 \$7206 \$7173 \$7147 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22940 \$153 \$7268 \$7173 \$7133 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22941 \$153 \$7032 \$5625 \$6677 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22942 \$153 \$7206 \$7463 \$7093 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22943 \$16 \$7147 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22944 \$16 \$7344 \$16 \$153 \$7093 VNB sky130_fd_sc_hd__inv_1
X$22945 \$16 \$7344 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22947 \$16 \$7130 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22948 \$16 \$7133 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22949 \$153 \$7092 \$7173 \$7131 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22950 \$153 \$7207 \$7173 \$7174 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22951 \$153 \$7207 \$7376 \$7093 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22952 \$153 \$7269 \$7639 \$7093 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22953 \$16 \$7174 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22956 \$153 \$7176 \$7240 \$7174 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22957 \$16 \$7131 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22958 \$153 \$7175 \$7208 \$7148 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22959 \$153 \$7176 \$7376 \$7148 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22961 \$153 \$7270 \$7240 \$7147 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22962 \$16 \$7174 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22963 \$16 \$7131 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22964 \$16 \$7130 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22968 \$153 \$7178 \$3199 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$22969 \$153 \$7271 \$7240 \$7133 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22970 \$16 \$7133 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22971 \$16 \$7178 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22973 \$16 \$7174 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22974 \$153 \$7179 \$3200 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$22976 \$16 \$7272 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22979 \$16 \$7709 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22980 \$16 \$7133 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22981 \$16 \$7147 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22982 \$153 \$7273 \$7241 \$7147 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22983 \$153 \$7177 \$7208 \$7097 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22984 \$153 \$7181 \$7241 \$7133 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22985 \$16 \$7179 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22988 \$153 \$7181 \$7180 \$7097 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22989 \$16 \$7174 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22990 \$153 \$7182 \$7242 \$7131 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22991 \$16 \$5636 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22992 \$153 \$7182 \$7208 \$7149 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$22993 \$153 \$7132 \$6619 \$5636 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22996 \$153 \$6923 \$6619 \$5963 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$22997 \$16 \$5609 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$22999 \$153 \$7132 \$5509 \$6639 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23000 \$153 \$7274 \$7243 \$7147 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23001 \$16 \$7147 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23002 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$23004 \$153 \$7183 \$7208 \$7392 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23005 \$153 \$7184 \$7243 \$7133 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23006 \$16 \$7133 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23007 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$23008 \$153 \$7184 \$7180 \$7392 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23009 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$23010 \$16 \$5609 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23012 \$16 \$7147 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23013 \$153 \$7050 \$5074 \$6633 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23015 \$153 \$7185 \$7244 \$7147 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23016 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$23018 \$153 \$7185 \$7463 \$6985 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23019 \$16 \$6985 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23021 \$16 \$7133 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23022 \$16 \$6985 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23023 \$153 \$7275 \$7244 \$7133 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23024 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$23025 \$16 \$7174 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23027 \$153 \$6975 \$7244 \$7174 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23028 \$153 \$7037 \$5806 \$6684 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23029 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$23030 \$153 \$6959 \$5074 \$6684 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23031 \$16 \$7174 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23032 \$16 \$7133 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23033 \$153 \$7209 \$7186 \$7174 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23036 \$153 \$7276 \$7186 \$7147 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23038 \$153 \$6897 \$5074 \$6565 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23039 \$16 \$7147 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23041 \$16 \$4954 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23042 \$153 \$5459 \$3142 \$4954 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23043 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$23044 \$16 \$5767 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23046 \$153 \$7134 \$6686 \$5767 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23047 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$23048 \$16 \$7147 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23049 \$153 \$7231 \$7245 \$7147 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23051 \$153 \$7134 \$5575 \$6561 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23052 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$23053 \$153 \$7038 \$5806 \$6561 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23054 \$16 \$7174 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23057 \$153 \$7232 \$7245 \$7174 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23058 \$153 \$6494 \$5509 \$6924 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23059 \$16 \$6924 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23060 \$153 \$6370 \$5484 \$6924 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23062 \$153 \$6395 \$5575 \$6924 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23066 \$153 \$7277 \$7187 \$7147 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23067 \$16 \$6924 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23068 \$16 \$6924 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23069 \$16 \$7147 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23070 \$153 \$6898 \$5938 \$6760 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23071 \$153 \$7210 \$7187 \$7131 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23072 \$16 \$4963 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23074 \$153 \$7052 \$5575 \$6760 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23076 \$16 \$7174 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23078 \$153 \$7211 \$7187 \$7174 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23079 \$153 \$7314 \$7187 \$7377 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23080 \$153 \$6748 \$5074 \$6457 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23082 \$153 \$7039 \$5509 \$6760 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23084 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$23085 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$23087 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$23088 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$23089 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$23090 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$23091 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$23093 \$153 \$7040 \$6859 \$6981 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23094 \$153 \$7018 \$6986 \$6783 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23095 \$153 \$7077 \$6930 \$7078 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23096 \$16 \$6783 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23097 \$16 \$6981 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23099 \$153 \$7019 \$6986 \$6860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23101 \$153 \$7018 \$6749 \$7078 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23102 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$23103 \$16 \$6860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23104 \$153 \$7100 \$6986 \$6792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23106 \$153 \$5663 \$5463 \$4579 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23108 \$16 \$4579 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23110 \$16 \$6792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23111 \$16 \$6987 \$16 \$153 \$6733 VNB sky130_fd_sc_hd__inv_1
X$23112 \$153 \$6927 \$6913 \$6709 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23113 \$153 \$6978 \$6781 \$7041 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23114 \$153 \$6781 \$6888 \$7101 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$23115 \$153 \$6978 \$6996 \$6709 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23117 \$16 \$6888 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23118 \$16 \$7041 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23119 \$16 \$7124 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23120 \$16 \$6987 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23121 \$16 \$6915 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23122 \$153 \$7054 \$7053 \$6979 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23123 \$153 \$6965 \$6781 \$6979 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23124 \$16 \$6988 \$16 \$153 \$6709 VNB sky130_fd_sc_hd__inv_1
X$23125 \$153 \$6859 \$6813 \$7102 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$23126 \$16 \$6979 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23128 \$153 \$6965 \$6995 \$6709 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23130 \$153 \$7103 \$6782 \$6981 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23131 \$153 \$7020 \$6782 \$7041 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23132 \$16 \$6981 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23133 \$153 \$6864 \$6719 \$6980 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23136 \$153 \$7020 \$6996 \$6980 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23138 \$16 \$6989 \$16 \$153 \$6980 VNB sky130_fd_sc_hd__inv_1
X$23139 \$153 \$6929 \$6995 \$6980 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23140 \$153 \$7103 \$6930 \$6980 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23141 \$153 \$6998 \$6751 \$7041 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23142 \$153 \$6997 \$6930 \$6815 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23144 \$153 \$6997 \$6751 \$6981 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23146 \$153 \$7104 \$6751 \$6979 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23147 \$153 \$6998 \$6996 \$6815 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23148 \$16 \$6979 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23149 \$16 \$7071 \$16 \$153 \$6815 VNB sky130_fd_sc_hd__inv_1
X$23150 \$16 \$6981 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23153 \$16 \$7071 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23154 \$153 \$6999 \$6752 \$7041 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23156 \$153 \$7021 \$6752 \$6979 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23157 \$16 \$7041 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23158 \$153 \$6999 \$6996 \$6692 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23159 \$153 \$7021 \$6995 \$6692 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23160 \$16 \$6979 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23162 \$153 \$7042 \$6752 \$6981 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23163 \$153 \$7042 \$6930 \$6692 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23164 \$153 \$7055 \$6908 \$7041 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23165 \$153 \$7022 \$6908 \$6907 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23166 \$16 \$6981 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23168 \$16 \$6909 \$16 \$153 \$6692 VNB sky130_fd_sc_hd__inv_1
X$23169 \$153 \$7055 \$6996 \$6914 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23170 \$16 \$7041 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23172 \$153 \$7105 \$6908 \$6979 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23173 \$16 \$6907 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23174 \$16 \$7000 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23175 \$16 \$6979 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23176 \$153 \$6934 \$6732 \$6914 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23178 \$153 \$7106 \$6785 \$6981 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23180 \$153 \$7022 \$6913 \$6914 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23181 \$153 \$7023 \$6785 \$6907 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23182 \$153 \$6785 \$7226 \$7056 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$23183 \$16 \$6935 \$16 \$153 \$6795 VNB sky130_fd_sc_hd__inv_1
X$23184 \$153 \$6902 \$6719 \$6795 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23186 \$16 \$6935 \$7158 \$7056 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$23187 \$16 \$7041 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23188 \$16 \$6907 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23189 \$153 \$7057 \$6786 \$6981 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23190 \$16 \$7226 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23191 \$153 \$6936 \$6913 \$6857 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23192 \$153 \$6886 \$6732 \$6857 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23193 \$153 \$7057 \$6930 \$6857 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23195 \$153 \$6966 \$6786 \$6792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23196 \$16 \$6910 \$7158 \$7107 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$23197 \$16 \$7072 \$16 \$153 \$6857 VNB sky130_fd_sc_hd__inv_1
X$23198 \$153 \$7001 \$6861 \$6979 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23200 \$153 \$6967 \$6861 \$6792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23202 \$16 \$6979 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23203 \$16 \$7072 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23204 \$153 \$6966 \$6719 \$6857 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23205 \$153 \$7108 \$6861 \$7041 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23206 \$153 \$6967 \$6719 \$6710 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23207 \$153 \$6796 \$6888 \$7024 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$23208 \$16 \$6988 \$6990 \$7024 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$23210 \$153 \$6968 \$6930 \$6710 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23211 \$153 \$7002 \$7073 \$6991 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23212 \$153 \$7001 \$6995 \$6710 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23213 \$153 \$6937 \$6913 \$6710 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23214 \$16 \$6988 \$16 \$153 \$6711 VNB sky130_fd_sc_hd__inv_1
X$23215 \$16 \$6991 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23216 \$153 \$7002 \$6992 \$6982 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23219 \$16 \$6988 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23220 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$23221 \$153 \$6969 \$6796 \$7060 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23222 \$153 \$7058 \$7073 \$6916 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23225 \$16 \$6916 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23226 \$153 \$7058 \$6867 \$6982 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23229 \$153 \$7192 \$6324 \$6982 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23231 \$16 \$6695 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23232 \$153 \$6938 \$6992 \$6711 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23233 \$153 \$7716 \$6787 \$7044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23235 \$153 \$7025 \$6787 \$6916 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23236 \$16 \$7044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23239 \$16 \$6987 \$16 \$153 \$6695 VNB sky130_fd_sc_hd__inv_1
X$23241 \$153 \$7079 \$6992 \$6695 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23242 \$153 \$6969 \$6324 \$6711 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23243 \$153 \$7059 \$7003 \$7043 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23244 \$16 \$6916 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23246 \$153 \$6889 \$7003 \$6713 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23247 \$153 \$7080 \$7003 \$7382 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23249 \$153 \$6970 \$6755 \$6991 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23250 \$153 \$6939 \$6867 \$6713 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23251 \$153 \$6651 \$6869 \$6862 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23252 \$153 \$6970 \$6992 \$6713 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23253 \$16 \$6991 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23254 \$16 \$6989 \$16 \$153 \$6652 VNB sky130_fd_sc_hd__inv_1
X$23256 \$153 \$7004 \$6869 \$6991 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23257 \$153 \$6800 \$6869 \$6771 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23258 \$153 \$7371 \$6869 \$7060 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23259 \$153 \$7004 \$6992 \$6652 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23262 \$16 \$6771 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23263 \$16 \$7071 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23264 \$16 \$7071 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23265 \$16 \$7071 \$16 \$153 \$6801 VNB sky130_fd_sc_hd__inv_1
X$23267 \$153 \$6871 \$6870 \$6771 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23268 \$16 \$7060 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23269 \$153 \$7061 \$6870 \$6991 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23271 \$153 \$6890 \$6906 \$6918 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23272 \$16 \$6991 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23275 \$153 \$7061 \$6992 \$6918 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23276 \$153 \$7005 \$7006 \$7043 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23277 \$16 \$7502 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23278 \$153 \$7007 \$6788 \$7044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23279 \$16 \$7399 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23281 \$16 \$6862 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23282 \$153 \$7007 \$7006 \$6801 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23284 \$153 \$7081 \$6324 \$6801 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23285 \$153 \$6891 \$6867 \$6801 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23286 \$16 \$7044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23287 \$153 \$6941 \$7003 \$6801 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23289 \$153 \$7009 \$6789 \$6991 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23291 \$153 \$7008 \$6324 \$6803 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23293 \$153 \$7009 \$6992 \$6803 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23294 \$16 \$6909 \$16 \$153 \$6803 VNB sky130_fd_sc_hd__inv_1
X$23296 \$153 \$7062 \$6789 \$7044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23297 \$153 \$6942 \$7003 \$6803 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23299 \$153 \$7010 \$7065 \$5932 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23300 \$153 \$7062 \$7006 \$6803 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23302 \$153 \$6804 \$6790 \$6862 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23303 \$16 \$7044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23304 \$153 \$7063 \$6790 \$7044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23305 \$16 \$6862 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23307 \$16 \$7044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23308 \$153 \$7063 \$7006 \$6805 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23310 \$16 \$6910 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23311 \$153 \$7026 \$6790 \$7060 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23313 \$153 \$7109 \$6790 \$6991 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23314 \$153 \$6831 \$6865 \$6805 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23315 \$16 \$6991 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23316 \$153 \$7011 \$6791 \$7060 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23317 \$16 \$7060 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23318 \$16 \$7072 \$16 \$153 \$6919 VNB sky130_fd_sc_hd__inv_1
X$23319 \$16 \$7072 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23322 \$16 \$7060 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23323 \$153 \$7011 \$6324 \$6919 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23324 \$16 \$6754 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23326 \$153 \$7012 \$6791 \$7044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23327 \$16 \$6991 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23328 \$153 \$7027 \$6791 \$6991 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23329 \$16 \$6797 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23333 \$153 \$7045 \$6791 \$6862 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23334 \$153 \$7027 \$6992 \$6919 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23335 \$153 \$6581 \$7013 \$7067 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23336 \$153 \$7012 \$7006 \$6919 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23338 \$153 \$7364 \$7366 \$5932 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23340 \$153 \$6135 \$7013 \$7129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23341 \$153 \$6583 \$7013 \$7029 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23342 \$16 \$7082 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23343 \$16 \$7129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23344 \$16 \$7029 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23345 \$153 \$7046 \$7014 \$7029 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23346 \$16 \$7029 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23347 \$16 \$5932 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23350 \$153 \$6945 \$5625 \$6556 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23353 \$16 \$7067 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23354 \$153 \$6971 \$6642 \$5702 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23355 \$153 \$7110 \$7014 \$7067 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23357 \$153 \$6971 \$5470 \$6556 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23358 \$16 \$5702 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23359 \$16 \$7082 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23360 \$16 \$5702 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23361 \$153 \$7145 \$6972 \$7082 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23362 \$153 \$7028 \$6972 \$7129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23363 \$16 \$7029 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23364 \$16 \$7129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23365 \$153 \$6946 \$5470 \$6616 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23369 \$16 \$7067 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23370 \$153 \$7167 \$6972 \$7067 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23371 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$23372 \$16 \$5605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23373 \$153 \$6973 \$6698 \$5605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23374 \$16 \$7082 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23375 \$153 \$7064 \$7074 \$7082 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23377 \$153 \$6973 \$5625 \$6616 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23378 \$153 \$7064 \$7065 \$7085 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23379 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$23381 \$153 \$6993 \$1677 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$23382 \$153 \$7083 \$7215 \$7085 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23385 \$153 \$7084 \$7066 \$7085 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23386 \$16 \$6993 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23388 \$16 \$5702 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23389 \$16 \$7067 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23390 \$153 \$6983 \$6643 \$5702 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23391 \$153 \$7111 \$7086 \$7067 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23393 \$153 \$7087 \$7086 \$7029 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23394 \$16 \$7029 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23395 \$16 \$6984 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23396 \$153 \$6983 \$5470 \$6714 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23398 \$153 \$6984 \$1678 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$23399 \$153 \$7087 \$7066 \$7112 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23400 \$16 \$7067 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23403 \$153 \$7088 \$7065 \$7112 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23405 \$153 \$6922 \$6511 \$5702 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23406 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$23407 \$153 \$7089 \$1544 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$23408 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$23411 \$153 \$7015 \$7066 \$7317 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23412 \$16 \$7089 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23413 \$16 \$7029 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23414 \$16 \$7067 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23415 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$23416 \$153 \$6644 \$7170 \$7067 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23417 \$16 \$5702 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23418 \$153 \$6974 \$6563 \$5702 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23421 \$16 \$7082 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23422 \$153 \$6775 \$5755 \$6533 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23423 \$153 \$7016 \$7171 \$7082 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23424 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$23425 \$153 \$7016 \$7065 \$7264 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23426 \$153 \$7075 \$1367 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$23427 \$16 \$5856 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23430 \$16 \$7129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23431 \$153 \$6839 \$5625 \$6560 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23432 \$153 \$7113 \$7090 \$7029 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23433 \$153 \$7047 \$7090 \$7129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23434 \$16 \$7075 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23437 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$23438 \$153 \$6950 \$5470 \$6560 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23439 \$16 \$7067 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23440 \$153 \$7114 \$7090 \$7067 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23441 \$153 \$7030 \$6742 \$5702 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23442 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$23443 \$16 \$7115 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23444 \$16 \$5702 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23446 \$153 \$7115 \$1673 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$23447 \$16 \$5400 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23448 \$16 \$5856 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23449 \$153 \$7031 \$6742 \$5856 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23450 \$153 \$7031 \$5795 \$6715 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23451 \$16 \$6269 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23452 \$16 \$6269 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23453 \$16 \$5173 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23454 \$16 \$5605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23456 \$153 \$7032 \$6703 \$5605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23457 \$153 \$7068 \$7065 \$6656 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23458 \$16 \$6656 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23460 \$153 \$7091 \$1516 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$23461 \$153 \$6953 \$5795 \$6677 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23463 \$16 \$7048 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23465 \$16 \$7386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23466 \$16 \$7033 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23467 \$16 \$5702 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23468 \$153 \$6954 \$5470 \$6677 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23469 \$16 \$1677 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23470 \$153 \$1677 \$5767 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$23471 \$16 \$7091 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23472 \$153 \$7092 \$7208 \$7093 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23473 \$16 \$7049 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23474 \$16 \$7033 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23475 \$153 \$6994 \$3243 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$23477 \$16 \$7033 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23478 \$153 \$7094 \$3439 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$23479 \$16 \$6994 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23480 \$16 \$1516 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23481 \$16 \$7094 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23483 \$16 \$7076 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23484 \$16 \$1678 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23485 \$16 \$7116 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23487 \$16 \$7069 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23488 \$153 \$1678 \$5963 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$23489 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$23490 \$153 \$7095 \$3508 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$23491 \$16 \$5609 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23492 \$16 \$4834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23494 \$16 \$5963 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23495 \$153 \$6896 \$5074 \$6657 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23497 \$16 \$7095 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23498 \$153 \$7096 \$7376 \$7097 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23500 \$153 \$6880 \$6681 \$5609 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23501 \$16 \$5609 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23502 \$16 \$7076 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23503 \$153 \$7034 \$3587 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$23504 \$16 \$6985 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23506 \$153 \$6956 \$5575 \$6682 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23507 \$153 \$7098 \$3720 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$23508 \$16 \$7034 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23510 \$16 \$5767 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23511 \$153 \$6975 \$7376 \$6985 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23512 \$153 \$7035 \$6619 \$5767 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23515 \$16 \$7098 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23516 \$16 \$5887 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23517 \$153 \$7035 \$5575 \$6639 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23518 \$153 \$6881 \$6619 \$5609 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23519 \$153 \$7099 \$3373 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$23522 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$23524 \$16 \$7099 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23525 \$16 \$5636 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23526 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$23527 \$153 \$7036 \$6631 \$5636 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23528 \$16 \$5767 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23529 \$153 \$7117 \$6631 \$5767 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23530 \$153 \$7050 \$6631 \$5609 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23532 \$153 \$7036 \$5509 \$6633 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23533 \$153 \$7117 \$5575 \$6633 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23535 \$153 \$7037 \$6640 \$5963 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23536 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$23537 \$16 \$5767 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23538 \$16 \$5636 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23539 \$153 \$7051 \$6640 \$5767 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23541 \$153 \$6976 \$6640 \$5636 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23542 \$153 \$7051 \$5575 \$6684 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23543 \$153 \$6976 \$5509 \$6684 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23544 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$23546 \$16 \$5636 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23547 \$16 \$5767 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23548 \$153 \$6977 \$6620 \$5636 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23550 \$153 \$7070 \$6620 \$5767 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23551 \$153 \$6977 \$5509 \$6565 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23552 \$153 \$7070 \$5575 \$6565 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23554 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$23555 \$16 \$5963 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23557 \$153 \$7038 \$6686 \$5963 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23559 \$16 \$5636 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23560 \$153 \$7017 \$6686 \$5636 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23561 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$23562 \$153 \$7017 \$5509 \$6561 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23563 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$23564 \$16 \$6924 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23568 \$16 \$5609 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23569 \$16 \$5636 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23570 \$153 \$6962 \$6688 \$5609 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23571 \$153 \$6925 \$6688 \$5636 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23573 \$16 \$5173 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23574 \$16 \$5963 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23576 \$153 \$6963 \$6688 \$5963 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23577 \$16 \$7131 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23578 \$16 \$5767 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23580 \$153 \$6926 \$6688 \$5767 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23581 \$16 \$5767 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23582 \$153 \$7118 \$6747 \$5963 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23583 \$153 \$7052 \$6747 \$5767 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23585 \$16 \$5963 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23586 \$16 \$7377 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23588 \$16 \$5636 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23589 \$16 \$5609 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23590 \$153 \$7119 \$6747 \$5609 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23591 \$153 \$7039 \$6747 \$5636 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23592 \$153 \$6690 \$5635 \$6457 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23593 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$23596 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$23597 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$23598 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$23599 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$23600 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$23601 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$23602 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$23603 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$23605 \$16 \$783 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23606 \$153 \$921 \$816 \$17 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23607 \$153 \$837 \$816 \$504 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23608 \$16 \$504 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23610 \$153 \$837 \$561 \$763 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23611 \$16 \$17 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23612 \$153 \$838 \$816 \$395 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23613 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$23614 \$16 \$710 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23615 \$153 \$838 \$394 \$763 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23616 \$16 \$395 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23618 \$16 \$710 \$503 \$780 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$23620 \$16 \$503 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23622 \$153 \$781 \$816 \$249 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23623 \$16 \$753 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23624 \$153 \$869 \$816 \$419 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23625 \$153 \$781 \$377 \$763 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23626 \$153 \$969 \$59 \$763 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23627 \$16 \$249 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23628 \$153 \$782 \$661 \$504 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23630 \$153 \$764 \$661 \$395 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23631 \$153 \$782 \$561 \$649 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23633 \$153 \$726 \$661 \$17 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23634 \$16 \$504 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23635 \$16 \$395 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23638 \$16 \$783 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23639 \$16 \$783 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23640 \$16 \$17 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23641 \$16 \$1291 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23642 \$153 \$870 \$661 \$184 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23643 \$153 \$784 \$661 \$58 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23644 \$153 \$784 \$30 \$649 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23645 \$16 \$184 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23646 \$16 \$537 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23649 \$153 \$870 \$59 \$649 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23650 \$16 \$58 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23651 \$16 \$754 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23652 \$16 \$582 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23653 \$16 \$582 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23655 \$16 \$541 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23656 \$153 \$839 \$755 \$58 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23657 \$153 \$922 \$755 \$249 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23659 \$153 \$923 \$755 \$419 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23660 \$16 \$249 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23662 \$153 \$554 \$394 \$96 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23664 \$153 \$681 \$817 \$504 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23665 \$153 \$839 \$30 \$903 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23667 \$16 \$249 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23669 \$153 \$840 \$817 \$395 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23670 \$153 \$924 \$817 \$17 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23671 \$153 \$785 \$349 \$639 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23672 \$16 \$17 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23674 \$16 \$58 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23676 \$153 \$871 \$664 \$263 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23677 \$16 \$395 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23679 \$153 \$787 \$664 \$58 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23680 \$16 \$263 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23681 \$153 \$872 \$664 \$395 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23682 \$153 \$787 \$30 \$765 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23683 \$153 \$786 \$377 \$765 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23685 \$16 \$899 \$16 \$153 \$765 VNB sky130_fd_sc_hd__inv_1
X$23686 \$16 \$395 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23688 \$16 \$899 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23689 \$153 \$887 \$561 \$651 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23690 \$16 \$1139 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23691 \$16 \$691 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23692 \$153 \$841 \$756 \$184 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23693 \$153 \$887 \$756 \$504 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23695 \$16 \$184 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23696 \$16 \$503 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23697 \$16 \$849 \$503 \$904 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$23698 \$16 \$842 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23699 \$16 \$849 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23700 \$16 \$504 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23701 \$153 \$788 \$756 \$249 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23703 \$153 \$873 \$756 \$419 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23704 \$153 \$788 \$377 \$651 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23707 \$16 \$849 \$16 \$153 \$651 VNB sky130_fd_sc_hd__inv_1
X$23708 \$16 \$419 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23709 \$16 \$249 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23711 \$153 \$843 \$583 \$395 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23712 \$153 \$874 \$583 \$263 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23713 \$16 \$395 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23714 \$153 \$843 \$394 \$766 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23716 \$16 \$504 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23718 \$153 \$844 \$583 \$504 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23719 \$16 \$263 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23720 \$16 \$652 \$715 \$818 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$23721 \$153 \$844 \$561 \$766 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23722 \$153 \$583 \$685 \$818 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$23723 \$153 \$888 \$349 \$173 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23726 \$153 \$506 \$584 \$729 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$23728 \$16 \$504 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23729 \$153 \$730 \$506 \$504 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23730 \$153 \$905 \$234 \$906 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23731 \$16 \$588 \$715 \$789 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$23732 \$153 \$433 \$506 \$395 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23733 \$16 \$395 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23735 \$153 \$889 \$506 \$17 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23736 \$153 \$889 \$102 \$432 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23737 \$16 \$280 \$555 \$790 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$23738 \$16 \$555 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23739 \$16 \$17 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23741 \$153 \$845 \$819 \$293 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23742 \$16 \$1037 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23743 \$16 \$1048 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23745 \$153 \$926 \$819 \$209 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23746 \$16 \$293 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23747 \$153 \$820 \$54 \$810 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23748 \$16 \$209 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23749 \$153 \$821 \$819 \$73 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23750 \$16 \$187 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23751 \$16 \$716 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23752 \$16 \$757 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23754 \$16 \$588 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23756 \$153 \$821 \$215 \$810 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23757 \$16 \$73 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23758 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$23759 \$153 \$927 \$819 \$212 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23760 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$23762 \$153 \$846 \$819 \$18 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23764 \$16 \$212 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23765 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$23766 \$16 \$18 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23767 \$153 \$907 \$104 \$810 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23768 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$23770 \$153 \$811 \$758 \$73 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23771 \$16 \$60 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23772 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$23774 \$153 \$928 \$758 \$60 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23777 \$153 \$811 \$215 \$767 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23778 \$16 \$60 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23780 \$153 \$847 \$758 \$187 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23781 \$153 \$768 \$758 \$18 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23783 \$16 \$582 \$16 \$153 \$105 VNB sky130_fd_sc_hd__inv_1
X$23785 \$153 \$847 \$54 \$767 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23786 \$16 \$187 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23787 \$16 \$18 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23788 \$153 \$587 \$753 \$822 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$23789 \$16 \$710 \$555 \$822 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$23790 \$16 \$555 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23791 \$153 \$812 \$587 \$73 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23792 \$16 \$753 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23793 \$16 \$710 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23794 \$16 \$507 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23795 \$16 \$582 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23798 \$153 \$812 \$215 \$600 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23799 \$16 \$73 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23800 \$16 \$187 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23802 \$16 \$18 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23803 \$16 \$710 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23804 \$153 \$875 \$823 \$18 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23805 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$23806 \$16 \$293 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23807 \$153 \$848 \$823 \$358 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23809 \$153 \$733 \$253 \$600 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23810 \$16 \$60 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23811 \$16 \$358 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23812 \$16 \$908 \$16 \$153 \$555 VNB sky130_fd_sc_hd__clkbuf_2
X$23813 \$153 \$572 \$347 \$600 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23814 \$153 \$690 \$1047 \$929 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$23815 \$153 \$734 \$346 \$600 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23816 \$153 \$876 \$900 \$209 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23818 \$16 \$555 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23819 \$16 \$1047 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23820 \$16 \$849 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23822 \$153 \$850 \$690 \$209 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23823 \$153 \$876 \$346 \$909 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23824 \$16 \$209 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23825 \$16 \$849 \$16 \$153 \$655 VNB sky130_fd_sc_hd__inv_1
X$23826 \$153 \$791 \$690 \$187 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23829 \$153 \$850 \$346 \$655 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23830 \$16 \$73 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23831 \$16 \$849 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23832 \$153 \$791 \$54 \$655 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23834 \$153 \$877 \$690 \$212 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23835 \$16 \$187 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23836 \$16 \$507 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23837 \$16 \$73 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23839 \$153 \$851 \$690 \$293 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23840 \$153 \$521 \$1659 \$930 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$23841 \$153 \$890 \$521 \$209 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23842 \$16 \$212 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23844 \$153 \$720 \$54 \$769 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23846 \$153 \$890 \$346 \$769 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23848 \$153 \$824 \$521 \$293 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23849 \$153 \$792 \$253 \$769 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23850 \$16 \$209 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23851 \$16 \$293 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23853 \$16 \$584 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23855 \$16 \$60 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23856 \$153 \$824 \$35 \$769 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23858 \$153 \$759 \$584 \$931 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$23859 \$16 \$652 \$946 \$793 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$23860 \$16 \$652 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23862 \$16 \$187 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23863 \$153 \$667 \$759 \$187 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23864 \$16 \$716 \$16 \$153 \$760 VNB sky130_fd_sc_hd__inv_1
X$23866 \$153 \$932 \$759 \$293 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23867 \$16 \$293 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23868 \$153 \$794 \$104 \$760 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23869 \$153 \$933 \$759 \$358 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23872 \$153 \$770 \$759 \$212 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23873 \$153 \$825 \$759 \$18 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23874 \$16 \$212 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23876 \$153 \$852 \$826 \$273 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23877 \$16 \$358 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23878 \$16 \$18 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23882 \$153 \$912 \$826 \$424 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23883 \$153 \$853 \$826 \$241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23884 \$153 \$878 \$826 \$145 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23885 \$16 \$79 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23886 \$16 \$273 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23889 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$23890 \$16 \$399 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23891 \$16 \$145 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23893 \$16 \$82 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23894 \$153 \$795 \$826 \$82 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23895 \$16 \$594 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23897 \$16 \$424 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23899 \$16 \$594 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23901 \$16 \$241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23903 \$16 \$273 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23904 \$153 \$855 \$854 \$241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23905 \$153 \$669 \$854 \$273 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23906 \$153 \$853 \$388 \$656 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23907 \$153 \$912 \$353 \$656 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23909 \$153 \$738 \$112 \$656 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23910 \$153 \$795 \$44 \$656 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23912 \$153 \$879 \$590 \$273 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23913 \$153 \$796 \$21 \$605 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23916 \$153 \$879 \$389 \$605 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23917 \$16 \$397 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23918 \$16 \$145 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23919 \$16 \$964 \$16 \$153 \$605 VNB sky130_fd_sc_hd__inv_1
X$23920 \$153 \$797 \$590 \$145 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23921 \$16 \$424 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23925 \$153 \$827 \$21 \$813 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23926 \$153 \$880 \$559 \$813 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23927 \$153 \$797 \$266 \$605 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23928 \$153 \$479 \$112 \$604 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23929 \$153 \$857 \$670 \$82 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23930 \$16 \$82 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23932 \$16 \$241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23934 \$153 \$936 \$670 \$241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23935 \$16 \$856 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23936 \$153 \$302 \$112 \$485 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23937 \$153 \$937 \$670 \$145 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23938 \$153 \$219 \$21 \$485 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23940 \$16 \$798 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23941 \$153 \$828 \$21 \$814 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23942 \$16 \$901 \$16 \$153 \$913 VNB sky130_fd_sc_hd__inv_1
X$23944 \$153 \$592 \$948 \$892 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$23946 \$16 \$424 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23947 \$153 \$799 \$592 \$424 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23948 \$16 \$829 \$268 \$892 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$23951 \$153 \$881 \$592 \$241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23953 \$153 \$858 \$592 \$273 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23954 \$16 \$241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23956 \$153 \$799 \$353 \$607 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23957 \$153 \$858 \$389 \$607 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23959 \$16 \$829 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23960 \$16 \$829 \$16 \$153 \$607 VNB sky130_fd_sc_hd__inv_1
X$23961 \$16 \$273 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23963 \$16 \$815 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23964 \$153 \$800 \$593 \$273 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23965 \$16 \$241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23966 \$153 \$744 \$593 \$241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23967 \$153 \$772 \$593 \$145 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23968 \$16 \$145 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23969 \$16 \$424 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23971 \$16 \$424 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23972 \$153 \$593 \$700 \$914 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$23974 \$16 \$815 \$16 \$153 \$771 VNB sky130_fd_sc_hd__inv_1
X$23975 \$153 \$801 \$830 \$82 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23976 \$16 \$82 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23977 \$153 \$859 \$353 \$611 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23979 \$153 \$859 \$830 \$424 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23980 \$153 \$938 \$353 \$915 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23982 \$153 \$830 \$895 \$894 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$23983 \$16 \$508 \$441 \$802 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$23985 \$16 \$241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23987 \$153 \$831 \$830 \$241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23990 \$153 \$831 \$388 \$611 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23991 \$153 \$916 \$21 \$915 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$23992 \$16 \$724 \$16 \$153 \$611 VNB sky130_fd_sc_hd__inv_1
X$23993 \$16 \$441 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23994 \$16 \$178 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23995 \$16 \$1303 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23996 \$153 \$804 \$761 \$178 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$23997 \$16 \$1120 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23998 \$16 \$1120 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$23999 \$16 \$508 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24000 \$16 \$895 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24001 \$16 \$446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24002 \$16 \$310 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24004 \$153 \$917 \$223 \$774 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24005 \$153 \$803 \$371 \$774 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24006 \$16 \$902 \$16 \$153 \$774 VNB sky130_fd_sc_hd__inv_1
X$24007 \$153 \$860 \$761 \$149 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24008 \$16 \$369 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24009 \$16 \$594 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24010 \$153 \$883 \$761 \$63 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24012 \$16 \$149 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24013 \$16 \$369 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24014 \$153 \$596 \$884 \$1016 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$24015 \$153 \$832 \$398 \$1087 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24016 \$16 \$63 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24017 \$16 \$178 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24018 \$153 \$861 \$596 \$178 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24019 \$153 \$939 \$703 \$774 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24022 \$153 \$896 \$371 \$658 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24023 \$153 \$861 \$549 \$658 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24024 \$153 \$885 \$596 \$63 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24025 \$153 \$860 \$398 \$774 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24026 \$16 \$63 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24028 \$153 \$885 \$57 \$658 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24029 \$16 \$509 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24031 \$153 \$702 \$223 \$658 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24032 \$16 \$901 \$428 \$940 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$24033 \$16 \$178 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24035 \$153 \$941 \$762 \$178 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24036 \$153 \$862 \$762 \$509 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24040 \$16 \$310 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24042 \$153 \$942 \$762 \$63 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24043 \$153 \$675 \$762 \$310 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24044 \$16 \$901 \$16 \$153 \$659 VNB sky130_fd_sc_hd__inv_1
X$24045 \$153 \$805 \$23 \$659 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24047 \$16 \$446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24048 \$16 \$178 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24049 \$153 \$886 \$706 \$178 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24051 \$153 \$833 \$57 \$775 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24052 \$153 \$806 \$23 \$775 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24053 \$153 \$886 \$549 \$775 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24054 \$153 \$660 \$427 \$63 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24055 \$16 \$63 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24056 \$16 \$798 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24057 \$16 \$428 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24060 \$16 \$815 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24061 \$16 \$509 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24062 \$153 \$863 \$706 \$509 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24063 \$16 \$309 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24064 \$153 \$834 \$706 \$309 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24066 \$16 \$829 \$428 \$864 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$24068 \$16 \$700 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24069 \$153 \$676 \$948 \$864 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$24071 \$153 \$834 \$703 \$775 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24072 \$16 \$178 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24073 \$153 \$807 \$676 \$178 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24074 \$153 \$863 \$371 \$775 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24075 \$16 \$615 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24076 \$16 \$815 \$615 \$897 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$24077 \$153 \$613 \$676 \$446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24079 \$153 \$943 \$700 \$897 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$24081 \$153 \$807 \$549 \$445 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24082 \$153 \$835 \$943 \$446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24084 \$16 \$829 \$16 \$153 \$445 VNB sky130_fd_sc_hd__inv_1
X$24087 \$153 \$835 \$393 \$776 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24088 \$153 \$777 \$676 \$509 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24089 \$153 \$865 \$836 \$509 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24090 \$153 \$866 \$57 \$779 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24091 \$153 \$866 \$836 \$63 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24093 \$153 \$778 \$836 \$309 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24094 \$16 \$724 \$615 \$867 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$24095 \$153 \$918 \$371 \$898 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24096 \$153 \$808 \$371 \$637 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24098 \$153 \$944 \$836 \$149 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24100 \$153 \$868 \$836 \$178 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24101 \$153 \$919 \$398 \$898 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24102 \$16 \$508 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24103 \$16 \$724 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24104 \$16 \$149 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24105 \$16 \$724 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24108 \$16 \$310 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24109 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$24110 \$153 \$920 \$223 \$898 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24111 \$153 \$809 \$23 \$779 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24112 \$153 \$725 \$393 \$779 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24113 \$153 \$868 \$549 \$779 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24114 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$24116 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$24117 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$24118 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$24119 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$24120 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$24121 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$24122 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$24123 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$24124 \$153 \$9600 \$9650 \$8950 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24125 \$153 \$9763 \$9650 \$8580 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24126 \$16 \$8950 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24127 \$16 \$8580 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24128 \$16 \$9129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24129 \$153 \$9734 \$8737 \$9728 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24130 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$24132 \$153 \$9601 \$9650 \$8828 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24134 \$153 \$9736 \$9650 \$8436 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24135 \$16 \$8828 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24136 \$16 \$8001 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24137 \$16 \$8114 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24138 \$16 \$9026 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24139 \$153 \$9799 \$8726 \$9728 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24140 \$16 \$8001 \$16 \$153 \$9392 VNB sky130_fd_sc_hd__inv_1
X$24142 \$153 \$9735 \$8209 \$9728 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24143 \$16 \$8436 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24144 \$16 \$8139 \$9547 \$9785 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$24145 \$153 \$9737 \$8457 \$9728 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24146 \$153 \$9831 \$8167 \$9785 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$24147 \$16 \$8001 \$9547 \$9715 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$24148 \$153 \$9331 \$9469 \$8436 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24149 \$16 \$8724 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24150 \$16 \$8167 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24152 \$153 \$10057 \$8209 \$9729 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24153 \$153 \$9800 \$8737 \$9729 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24154 \$153 \$9716 \$8457 \$9729 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24155 \$153 \$9832 \$8503 \$9764 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$24156 \$16 \$8423 \$9547 \$9764 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$24157 \$16 \$8436 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24160 \$153 \$9394 \$9469 \$9026 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24161 \$16 \$8724 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24162 \$16 \$8503 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24164 \$16 \$8423 \$16 \$153 \$9583 VNB sky130_fd_sc_hd__inv_1
X$24165 \$153 \$9680 \$9543 \$8828 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24166 \$16 \$9026 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24167 \$16 \$8724 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24168 \$16 \$8715 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24169 \$153 \$9717 \$9543 \$8715 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24171 \$16 \$8828 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24172 \$16 \$8423 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24174 \$153 \$9833 \$8912 \$9449 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24175 \$153 \$9717 \$8638 \$9449 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24176 \$16 \$8950 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24178 \$153 \$9681 \$9543 \$8436 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24179 \$153 \$9738 \$8737 \$9583 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24181 \$153 \$9765 \$8297 \$9739 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$24182 \$16 \$8144 \$9547 \$9739 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$24183 \$16 \$8436 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24184 \$153 \$9801 \$9765 \$9129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24186 \$153 \$9766 \$9765 \$8724 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24189 \$153 \$9801 \$8737 \$9740 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24190 \$16 \$8144 \$16 \$153 \$9740 VNB sky130_fd_sc_hd__inv_1
X$24191 \$16 \$8724 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24193 \$153 \$9767 \$9459 \$8724 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24194 \$16 \$9129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24195 \$153 \$9802 \$9793 \$8724 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24196 \$16 \$8724 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24199 \$153 \$9638 \$8209 \$9321 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24201 \$16 \$8118 \$9260 \$9803 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$24202 \$153 \$9595 \$9606 \$8436 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24203 \$153 \$9768 \$9606 \$9026 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24204 \$16 \$8436 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24205 \$16 \$8118 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24206 \$153 \$9768 \$8726 \$9585 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24207 \$16 \$8118 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24209 \$16 \$8025 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24210 \$16 \$8177 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24211 \$16 \$8177 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24212 \$16 \$9026 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24213 \$16 \$9129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24215 \$153 \$9718 \$9606 \$8828 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24216 \$153 \$9786 \$9606 \$9129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24217 \$153 \$9786 \$8737 \$9585 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24218 \$16 \$8828 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24221 \$153 \$9718 \$8885 \$9585 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24222 \$16 \$8828 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24223 \$16 \$8177 \$9260 \$9804 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$24224 \$153 \$9565 \$8457 \$9585 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24225 \$153 \$9880 \$8169 \$9804 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$24226 \$16 \$7535 \$9260 \$9607 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$24228 \$153 \$9769 \$9673 \$8580 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24229 \$16 \$8580 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24231 \$153 \$9838 \$8061 \$9837 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$24232 \$153 \$9741 \$9673 \$8436 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24233 \$153 \$9805 \$8737 \$9867 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24234 \$16 \$9129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24235 \$16 \$8724 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24237 \$16 \$8724 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24238 \$153 \$9683 \$8638 \$9567 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24240 \$153 \$9806 \$8457 \$9867 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24242 \$16 \$10042 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24243 \$153 \$9769 \$8194 \$9567 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24244 \$16 \$8885 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24246 \$153 \$9684 \$9673 \$8950 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24247 \$16 \$8125 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24248 \$16 \$8457 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24249 \$16 \$8912 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24250 \$16 \$8194 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24252 \$16 \$9129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24253 \$16 \$8950 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24254 \$153 \$9770 \$9673 \$9129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24255 \$16 \$8209 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24256 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24257 \$153 \$9807 \$8340 \$8457 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24258 \$153 \$9655 \$8726 \$9567 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24259 \$153 \$9808 \$9787 \$8886 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24262 \$153 \$9548 \$9609 \$8886 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24263 \$153 \$9787 \$7884 \$9771 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$24264 \$16 \$8001 \$9371 \$9771 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$24266 \$153 \$9719 \$9609 \$8647 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24267 \$16 \$8886 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24269 \$153 \$9610 \$9787 \$8647 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24270 \$153 \$9719 \$8614 \$9533 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24272 \$153 \$9612 \$9609 \$8728 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24273 \$16 \$8647 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24274 \$16 \$8647 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24275 \$16 \$8139 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24276 \$16 \$8728 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24278 \$153 \$9742 \$9609 \$8556 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24279 \$153 \$9534 \$9787 \$8686 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24280 \$153 \$9742 \$8610 \$9533 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24281 \$16 \$8139 \$9371 \$9788 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$24282 \$16 \$8556 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24283 \$16 \$8686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24284 \$153 \$9462 \$9481 \$8816 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24286 \$153 \$9743 \$9794 \$8728 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24287 \$153 \$9743 \$8818 \$9902 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24288 \$153 \$9794 \$8167 \$9788 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$24289 \$16 \$8816 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24290 \$16 \$8728 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24292 \$16 \$8271 \$9371 \$9772 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$24293 \$153 \$9730 \$9795 \$8728 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24295 \$153 \$9730 \$8818 \$9720 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24296 \$153 \$9618 \$9484 \$8728 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24297 \$153 \$9840 \$8614 \$9720 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24300 \$16 \$8271 \$16 \$153 \$9720 VNB sky130_fd_sc_hd__inv_1
X$24301 \$16 \$8728 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24302 \$153 \$9809 \$9796 \$8728 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24303 \$16 \$8728 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24305 \$153 \$9619 \$9484 \$8886 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24306 \$16 \$8728 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24307 \$16 \$8271 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24309 \$16 \$8886 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24310 \$16 \$8169 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24312 \$153 \$9811 \$8169 \$9810 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$24314 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$24315 \$16 \$8177 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24316 \$153 \$9773 \$9487 \$8647 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24317 \$153 \$9596 \$9811 \$8728 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24318 \$16 \$8647 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24319 \$153 \$9744 \$8727 \$9586 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24321 \$153 \$9812 \$8610 \$9586 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24322 \$153 \$9721 \$9487 \$8890 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24323 \$16 \$8125 \$9400 \$9813 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$24324 \$153 \$9884 \$8061 \$9813 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$24325 \$16 \$8890 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24326 \$16 \$8061 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24327 \$16 \$8125 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24330 \$153 \$9814 \$8610 \$9815 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24331 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$24333 \$153 \$9640 \$8818 \$9421 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24334 \$153 \$9687 \$8804 \$9488 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24335 \$153 \$9688 \$9463 \$8686 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24337 \$153 \$9789 \$8818 \$9815 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24339 \$153 \$9846 \$8025 \$9844 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$24340 \$16 \$8686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24341 \$16 \$8125 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24342 \$16 \$8025 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24343 \$153 \$9689 \$9403 \$8898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24344 \$153 \$9816 \$9403 \$8816 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24345 \$16 \$8898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24347 \$16 \$8890 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24349 \$16 \$8816 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24350 \$153 \$9847 \$9403 \$8886 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24351 \$153 \$9774 \$9403 \$8728 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24352 \$153 \$9816 \$8804 \$9452 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24353 \$16 \$8886 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24354 \$16 \$8686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24355 \$153 \$9745 \$9660 \$8686 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24357 \$153 \$9848 \$9660 \$8886 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24358 \$153 \$9774 \$8818 \$9452 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24359 \$16 \$8816 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24360 \$16 \$7535 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24361 \$16 \$7535 \$16 \$153 \$9746 VNB sky130_fd_sc_hd__inv_1
X$24362 \$16 \$8728 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24363 \$153 \$9748 \$9660 \$8728 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24364 \$16 \$8556 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24365 \$16 \$8647 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24367 \$153 \$9775 \$9660 \$8647 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24368 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24369 \$153 \$9569 \$8340 \$10501 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24370 \$16 \$9747 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24371 \$153 \$9747 \$9275 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$24373 \$153 \$8670 \$8936 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$24374 \$16 \$9138 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24375 \$153 \$9722 \$9732 \$8807 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24376 \$153 \$9138 \$9253 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$24378 \$153 \$8516 \$9045 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$24379 \$153 \$9775 \$8614 \$9746 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24380 \$153 \$9748 \$8818 \$9746 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24381 \$16 \$9045 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24382 \$16 \$9253 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24383 \$16 \$16 \$153 VNB sky130_fd_sc_hd__conb_1
X$24386 \$153 \$153 \$9047 \$9625 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24387 \$153 \$153 \$9174 \$9625 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24388 \$153 \$153 \$8842 \$9625 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24390 \$153 \$9732 \$7839 \$9849 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$24391 \$153 \$153 \$8917 \$9625 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24392 \$153 \$9662 \$9693 \$8807 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24394 \$153 \$9692 \$9693 \$9045 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24395 \$153 \$9850 \$9252 \$9587 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24396 \$16 \$8220 \$9518 \$9723 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$24398 \$16 \$8936 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24399 \$153 \$9626 \$9693 \$8936 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24400 \$16 \$9253 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24401 \$16 \$9031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24403 \$153 \$9454 \$9693 \$9031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24404 \$16 \$8673 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24405 \$153 \$9749 \$9278 \$9587 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24407 \$153 \$9750 \$9674 \$8936 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24408 \$16 \$8936 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24410 \$16 \$8044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24411 \$16 \$7904 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24413 \$16 \$9188 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24414 \$16 \$8807 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24415 \$153 \$9750 \$8842 \$9695 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24416 \$16 \$8250 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24417 \$16 \$9188 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24418 \$16 \$8044 \$16 \$153 \$9695 VNB sky130_fd_sc_hd__inv_1
X$24419 \$153 \$9627 \$9674 \$9188 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24420 \$16 \$9045 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24421 \$153 \$9553 \$9674 \$8807 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24423 \$153 \$9851 \$9133 \$9695 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24425 \$16 \$7904 \$9518 \$9628 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$24427 \$153 \$9696 \$9544 \$9188 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24428 \$16 \$9214 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24429 \$153 \$9818 \$9047 \$9465 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24430 \$153 \$9797 \$9544 \$9275 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24431 \$16 \$8936 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24433 \$16 \$9031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24434 \$16 \$9188 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24435 \$16 \$9188 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24436 \$153 \$9751 \$9252 \$9465 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24437 \$153 \$9797 \$9278 \$9465 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24439 \$153 \$9724 \$9466 \$9188 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24440 \$16 \$8936 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24441 \$153 \$9853 \$9278 \$9642 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24443 \$153 \$9852 \$9752 \$8936 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24444 \$153 \$9776 \$9752 \$9031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24446 \$153 \$10022 \$8702 \$9854 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$24448 \$16 \$8316 \$9733 \$9697 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$24449 \$16 \$9253 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24451 \$153 \$9753 \$9047 \$9642 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24452 \$16 \$9253 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24453 \$153 \$9819 \$9752 \$9253 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24454 \$16 \$9275 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24455 \$153 \$9777 \$9433 \$9253 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24456 \$16 \$8702 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24457 \$16 \$8453 \$9733 \$9754 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$24458 \$16 \$8316 \$16 \$153 \$9642 VNB sky130_fd_sc_hd__inv_1
X$24460 \$153 \$9777 \$9252 \$9521 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24461 \$16 \$8453 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24463 \$153 \$9755 \$8732 \$9754 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$24464 \$16 \$8732 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24465 \$16 \$9031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24466 \$153 \$9820 \$9755 \$9031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24467 \$153 \$9756 \$8676 \$9725 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24469 \$153 \$9631 \$9408 \$9031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24470 \$153 \$9820 \$9133 \$9725 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24471 \$16 \$8936 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24472 \$153 \$9821 \$9755 \$8936 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24473 \$153 \$9757 \$9174 \$9642 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24474 \$16 \$8704 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24475 \$16 \$8453 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24477 \$16 \$8453 \$16 \$153 \$9725 VNB sky130_fd_sc_hd__inv_1
X$24478 \$153 \$9821 \$8842 \$9725 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24479 \$153 \$9667 \$8917 \$9409 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24480 \$153 \$9855 \$9174 \$9725 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24481 \$153 \$9758 \$8473 \$9698 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$24483 \$153 \$9822 \$8917 \$9823 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24486 \$153 \$9731 \$9524 \$9214 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24487 \$153 \$9778 \$9758 \$9045 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24488 \$153 \$9731 \$9047 \$9555 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24489 \$153 \$9778 \$9174 \$9823 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24490 \$16 \$9031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24491 \$16 \$9031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24493 \$153 \$9699 \$9524 \$9031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24495 \$153 \$9790 \$9758 \$9275 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24497 \$153 \$9577 \$8842 \$9555 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24498 \$16 \$8265 \$16 \$153 \$9823 VNB sky130_fd_sc_hd__inv_1
X$24499 \$16 \$9275 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24500 \$16 \$8265 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24501 \$153 \$153 \$9059 \$9701 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24502 \$16 \$8359 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24505 \$16 \$8473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24507 \$153 \$153 \$8965 \$9701 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24508 \$153 \$153 \$8996 \$9701 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24509 \$16 \$8719 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24510 \$16 \$16 \$153 VNB sky130_fd_sc_hd__conb_1
X$24511 \$153 \$153 \$9103 \$9701 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24513 \$153 \$153 \$8977 \$9701 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24514 \$16 \$8996 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24515 \$16 \$8187 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24516 \$153 \$153 \$9256 \$9701 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24518 \$153 \$153 \$9122 \$9701 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24519 \$16 \$8673 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24520 \$153 \$9779 \$9702 \$9134 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24521 \$153 \$9824 \$9702 \$9035 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24523 \$16 \$9035 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24524 \$16 \$8927 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24526 \$153 \$9824 \$8977 \$9759 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24527 \$16 \$8187 \$16 \$153 \$9759 VNB sky130_fd_sc_hd__inv_1
X$24528 \$16 \$9134 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24530 \$153 \$9780 \$9702 \$8879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24531 \$153 \$9857 \$9256 \$9759 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24532 \$16 \$9154 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24533 \$153 \$9780 \$8923 \$9759 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24534 \$16 \$8879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24536 \$153 \$9760 \$9702 \$9034 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24538 \$153 \$9825 \$9702 \$9154 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24539 \$153 \$9671 \$8965 \$9759 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24540 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$24541 \$16 \$9035 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24542 \$153 \$9826 \$9676 \$9035 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24543 \$16 \$9034 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24545 \$16 \$9134 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24547 \$153 \$9559 \$9676 \$9134 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24548 \$153 \$9760 \$9059 \$9759 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24549 \$153 \$9703 \$9676 \$8844 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24550 \$153 \$9826 \$8977 \$9560 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24553 \$16 \$9035 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24554 \$153 \$9827 \$9103 \$9560 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24555 \$16 \$8844 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24556 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$24557 \$16 \$9134 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24559 \$153 \$9635 \$9677 \$9134 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24560 \$153 \$9828 \$9677 \$9035 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24562 \$153 \$9828 \$8977 \$9592 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24564 \$16 \$9034 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24565 \$153 \$9704 \$9256 \$9592 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24567 \$16 \$9154 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24568 \$153 \$9829 \$9677 \$9154 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24570 \$153 \$9761 \$9677 \$9034 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24572 \$153 \$9829 \$9103 \$9592 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24573 \$153 \$9705 \$8965 \$9592 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24574 \$153 \$9726 \$8705 \$9762 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$24575 \$16 \$9035 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24576 \$16 \$8165 \$9562 \$9762 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$24577 \$153 \$9859 \$9726 \$9035 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24579 \$16 \$8165 \$16 \$153 \$9708 VNB sky130_fd_sc_hd__inv_1
X$24581 \$153 \$9761 \$9059 \$9592 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24582 \$16 \$8165 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24583 \$16 \$9798 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24584 \$16 \$8285 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24586 \$16 \$8893 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24587 \$16 \$8844 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24588 \$153 \$9727 \$9726 \$8844 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24589 \$153 \$9707 \$9726 \$8893 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24592 \$153 \$9727 \$8965 \$9708 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24593 \$16 \$9034 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24594 \$16 \$8732 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24595 \$153 \$9860 \$8732 \$9791 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$24597 \$153 \$9678 \$8285 \$9643 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$24598 \$16 \$8453 \$9562 \$9791 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$24599 \$153 \$9862 \$9678 \$9035 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24600 \$16 \$9035 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24603 \$153 \$10176 \$9678 \$8927 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24604 \$16 \$8453 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24606 \$16 \$8316 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24607 \$16 \$8316 \$16 \$153 \$10222 VNB sky130_fd_sc_hd__inv_1
X$24609 \$16 \$8893 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24610 \$153 \$8551 \$7462 \$8266 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24612 \$153 \$9781 \$9678 \$8893 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24614 \$16 \$8266 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24615 \$16 \$8359 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24617 \$16 \$9134 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24618 \$153 \$9782 \$9678 \$9134 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24620 \$153 \$8269 \$7376 \$8266 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24621 \$153 \$9792 \$8473 \$9711 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$24622 \$16 \$8266 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24623 \$16 \$8359 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24625 \$16 \$8473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24626 \$16 \$9134 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24627 \$16 \$8266 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24628 \$153 \$9783 \$9792 \$9134 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24629 \$16 \$8879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24630 \$153 \$9863 \$9792 \$8879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24631 \$16 \$9154 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24632 \$153 \$8778 \$7639 \$8777 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24633 \$16 \$8265 \$16 \$153 \$10510 VNB sky130_fd_sc_hd__inv_1
X$24634 \$16 \$9034 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24636 \$153 \$9830 \$9581 \$9034 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24637 \$153 \$9784 \$9581 \$9154 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24638 \$153 \$11054 \$9792 \$9035 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24639 \$153 \$9648 \$9059 \$9366 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24641 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$24643 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$24644 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$24645 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$24646 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$24647 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$24648 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$24649 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$24650 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$24652 \$153 \$231 \$234 \$88 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24655 \$153 \$231 \$64 \$263 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24656 \$153 \$202 \$64 \$58 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24658 \$153 \$202 \$30 \$88 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24659 \$16 \$263 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24660 \$16 \$58 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24661 \$16 \$264 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24662 \$16 \$395 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24665 \$16 \$264 \$16 \$153 \$88 VNB sky130_fd_sc_hd__inv_1
X$24666 \$153 \$246 \$64 \$249 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24667 \$153 \$246 \$377 \$88 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24668 \$153 \$127 \$59 \$88 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24669 \$153 \$90 \$65 \$58 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24670 \$16 \$249 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24671 \$16 \$419 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24673 \$16 \$263 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24676 \$153 \$247 \$65 \$249 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24677 \$153 \$203 \$65 \$184 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24678 \$16 \$249 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24679 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$24680 \$16 \$184 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24681 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$24682 \$153 \$92 \$182 \$249 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24684 \$153 \$91 \$182 \$184 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24685 \$153 \$278 \$234 \$89 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24686 \$16 \$184 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24687 \$153 \$93 \$182 \$17 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24688 \$16 \$249 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24689 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$24692 \$153 \$205 \$30 \$94 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24693 \$153 \$205 \$182 \$58 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24694 \$16 \$279 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24695 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$24696 \$153 \$95 \$66 \$58 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24697 \$16 \$58 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24698 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$24700 \$153 \$206 \$66 \$184 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24701 \$153 \$128 \$102 \$96 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24702 \$16 \$58 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24703 \$16 \$279 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24704 \$16 \$184 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24705 \$16 \$280 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24706 \$153 \$97 \$67 \$17 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24707 \$153 \$248 \$377 \$270 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24709 \$153 \$248 \$67 \$249 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24710 \$153 \$207 \$67 \$184 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24711 \$153 \$207 \$59 \$270 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24712 \$16 \$184 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24713 \$16 \$17 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24714 \$16 \$184 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24716 \$153 \$281 \$68 \$249 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24718 \$153 \$154 \$68 \$58 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24719 \$153 \$154 \$30 \$98 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24720 \$153 \$131 \$102 \$98 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24721 \$16 \$249 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24722 \$16 \$58 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24723 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$24725 \$153 \$155 \$190 \$58 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24727 \$153 \$99 \$190 \$184 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24729 \$153 \$155 \$30 \$100 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24730 \$153 \$191 \$190 \$263 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24731 \$16 \$184 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24733 \$153 \$191 \$234 \$100 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24734 \$16 \$263 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24736 \$153 \$282 \$69 \$249 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24737 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$24739 \$153 \$156 \$69 \$58 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24740 \$16 \$249 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24741 \$16 \$58 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24743 \$153 \$250 \$69 \$263 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24744 \$153 \$156 \$30 \$101 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24745 \$153 \$183 \$59 \$101 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24747 \$153 \$251 \$70 \$249 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24748 \$16 \$263 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24750 \$16 \$263 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24753 \$153 \$132 \$102 \$172 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24754 \$153 \$251 \$377 \$172 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24755 \$153 \$103 \$70 \$184 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24756 \$153 \$283 \$349 \$172 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24757 \$16 \$249 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24759 \$16 \$395 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24760 \$16 \$184 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24762 \$16 \$249 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24763 \$153 \$284 \$71 \$263 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24764 \$153 \$157 \$71 \$249 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24765 \$16 \$263 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24766 \$153 \$157 \$377 \$173 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24767 \$16 \$58 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24768 \$16 \$264 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24769 \$16 \$184 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24770 \$153 \$285 \$71 \$184 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24773 \$153 \$158 \$71 \$17 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24774 \$16 \$555 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24775 \$16 \$264 \$555 \$286 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$24776 \$153 \$158 \$102 \$173 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24777 \$153 \$320 \$54 \$271 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24779 \$153 \$159 \$72 \$209 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24781 \$153 \$287 \$72 \$293 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24782 \$153 \$159 \$346 \$174 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24783 \$16 \$187 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24784 \$16 \$293 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24785 \$16 \$588 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24786 \$153 \$252 \$72 \$358 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24787 \$16 \$209 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24788 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$24790 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$24791 \$153 \$133 \$215 \$174 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24792 \$153 \$252 \$253 \$174 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24793 \$16 \$358 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24794 \$153 \$160 \$72 \$18 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24795 \$153 \$321 \$215 \$271 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24797 \$153 \$288 \$420 \$18 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24798 \$16 \$18 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24799 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$24800 \$16 \$18 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24802 \$153 \$236 \$74 \$18 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24804 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$24806 \$16 \$18 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24807 \$153 \$134 \$104 \$175 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24808 \$153 \$52 \$185 \$73 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24809 \$153 \$135 \$215 \$175 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24810 \$153 \$161 \$185 \$60 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24811 \$16 \$73 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24812 \$16 \$507 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24814 \$153 \$289 \$185 \$209 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24815 \$153 \$161 \$104 \$105 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24816 \$16 \$209 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24817 \$16 \$293 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24818 \$16 \$60 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24819 \$153 \$272 \$192 \$73 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24820 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$24822 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$24823 \$153 \$210 \$192 \$60 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24824 \$153 \$290 \$192 \$187 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24825 \$153 \$211 \$192 \$18 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24826 \$16 \$60 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24827 \$16 \$73 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24829 \$153 \$291 \$24 \$212 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24830 \$16 \$212 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24831 \$153 \$213 \$24 \$73 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24832 \$153 \$292 \$24 \$209 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24835 \$153 \$137 \$104 \$325 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24836 \$153 \$213 \$215 \$325 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24837 \$16 \$209 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24838 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$24839 \$153 \$272 \$215 \$186 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24840 \$153 \$163 \$53 \$60 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24841 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$24842 \$16 \$293 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24844 \$16 \$212 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24845 \$153 \$163 \$104 \$176 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24846 \$153 \$138 \$215 \$176 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24847 \$153 \$19 \$193 \$187 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24848 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$24850 \$16 \$187 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24851 \$153 \$238 \$193 \$212 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24853 \$16 \$187 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24854 \$153 \$238 \$347 \$20 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24855 \$153 \$107 \$193 \$18 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24856 \$153 \$195 \$193 \$73 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24857 \$16 \$209 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24858 \$16 \$212 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24859 \$16 \$18 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24860 \$16 \$73 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24864 \$153 \$214 \$194 \$209 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24865 \$16 \$293 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24866 \$153 \$164 \$194 \$18 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24867 \$153 \$195 \$215 \$20 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24868 \$16 \$209 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24869 \$16 \$18 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24870 \$153 \$239 \$194 \$187 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24873 \$153 \$216 \$194 \$60 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24874 \$153 \$216 \$104 \$188 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24875 \$16 \$60 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24876 \$16 \$73 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24878 \$16 \$187 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24879 \$153 \$217 \$75 \$187 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24880 \$16 \$187 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24881 \$16 \$358 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24882 \$16 \$293 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24884 \$153 \$294 \$75 \$293 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24885 \$153 \$239 \$54 \$188 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24886 \$153 \$240 \$75 \$209 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24889 \$153 \$108 \$75 \$18 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24890 \$153 \$295 \$75 \$212 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24891 \$153 \$240 \$346 \$329 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24892 \$16 \$212 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24893 \$16 \$358 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24895 \$16 \$18 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24896 \$16 \$273 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24899 \$153 \$296 \$76 \$273 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24900 \$153 \$196 \$76 \$145 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24902 \$153 \$196 \$266 \$352 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24904 \$16 \$82 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24905 \$153 \$109 \$76 \$82 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24907 \$153 \$297 \$76 \$241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24908 \$153 \$218 \$559 \$352 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24909 \$16 \$241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24910 \$16 \$145 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24912 \$16 \$273 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24914 \$16 \$82 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24917 \$153 \$299 \$61 \$273 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24918 \$153 \$110 \$61 \$82 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24919 \$153 \$140 \$112 \$352 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24920 \$16 \$397 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24921 \$16 \$595 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24922 \$16 \$265 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24923 \$16 \$424 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24924 \$153 \$254 \$61 \$424 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24927 \$153 \$254 \$353 \$111 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24928 \$153 \$165 \$559 \$111 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24929 \$16 \$265 \$16 \$153 \$111 VNB sky130_fd_sc_hd__inv_1
X$24931 \$16 \$241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24932 \$153 \$166 \$77 \$82 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24934 \$153 \$255 \$77 \$145 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24935 \$153 \$166 \$44 \$113 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24936 \$153 \$255 \$266 \$113 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24937 \$16 \$79 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24938 \$16 \$145 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24940 \$16 \$423 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24941 \$16 \$265 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24942 \$153 \$143 \$21 \$113 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24943 \$153 \$300 \$78 \$145 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24946 \$153 \$301 \$78 \$79 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24947 \$153 \$197 \$44 \$115 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24948 \$153 \$167 \$21 \$115 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24949 \$16 \$79 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24951 \$16 \$82 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24952 \$153 \$303 \$189 \$82 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24954 \$16 \$151 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24956 \$16 \$151 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24957 \$16 \$79 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24958 \$153 \$302 \$189 \$79 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24959 \$16 \$268 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24961 \$153 \$198 \$21 \$177 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24962 \$16 \$82 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24964 \$153 \$256 \$267 \$82 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24965 \$153 \$144 \$559 \$177 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24966 \$153 \$274 \$266 \$177 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24967 \$153 \$256 \$44 \$177 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24968 \$16 \$273 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24969 \$153 \$304 \$267 \$273 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24971 \$16 \$80 \$268 \$410 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$24973 \$16 \$82 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24975 \$153 \$220 \$559 \$117 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24976 \$153 \$119 \$81 \$145 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24978 \$16 \$268 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24980 \$153 \$305 \$353 \$117 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24981 \$16 \$1456 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24984 \$16 \$273 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24985 \$153 \$336 \$388 \$117 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24986 \$153 \$221 \$62 \$273 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24987 \$16 \$424 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24988 \$16 \$306 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24990 \$16 \$258 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24991 \$153 \$221 \$389 \$120 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24993 \$16 \$79 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$24994 \$153 \$222 \$62 \$79 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$24997 \$153 \$147 \$559 \$120 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$24998 \$16 \$276 \$16 \$153 \$120 VNB sky130_fd_sc_hd__inv_1
X$24999 \$153 \$168 \$62 \$145 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25000 \$153 \$257 \$62 \$241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25002 \$153 \$257 \$388 \$120 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25003 \$153 \$168 \$266 \$120 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25005 \$153 \$244 \$57 \$258 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25007 \$16 \$310 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25008 \$153 \$169 \$83 \$310 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25009 \$153 \$22 \$223 \$258 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25011 \$153 \$224 \$549 \$121 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25012 \$153 \$224 \$83 \$178 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25013 \$153 \$259 \$83 \$446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25014 \$153 \$169 \$223 \$121 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25015 \$153 \$259 \$393 \$121 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25018 \$153 \$225 \$83 \$149 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25020 \$153 \$243 \$84 \$149 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25022 \$16 \$63 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25023 \$16 \$178 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25026 \$153 \$307 \$84 \$178 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25027 \$153 \$244 \$84 \$63 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25028 \$16 \$428 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25030 \$16 \$178 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25031 \$16 \$310 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25032 \$153 \$308 \$85 \$178 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25033 \$16 \$149 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25035 \$16 \$149 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25037 \$153 \$123 \$85 \$149 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25039 \$16 \$309 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25040 \$153 \$199 \$85 \$309 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25041 \$16 \$428 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25042 \$16 \$354 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25043 \$153 \$199 \$703 \$122 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25046 \$153 \$148 \$23 \$122 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25047 \$153 \$275 \$703 \$124 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25048 \$153 \$260 \$227 \$310 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25049 \$16 \$265 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25050 \$153 \$260 \$223 \$124 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25052 \$16 \$354 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25053 \$16 \$149 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25054 \$153 \$200 \$227 \$149 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25056 \$153 \$311 \$227 \$178 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25057 \$16 \$178 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25058 \$16 \$151 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25060 \$16 \$591 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25061 \$16 \$178 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25062 \$153 \$312 \$86 \$178 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25063 \$153 \$228 \$86 \$310 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25065 \$16 \$310 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25066 \$16 \$309 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25068 \$153 \$200 \$398 \$124 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25069 \$153 \$1180 \$86 \$309 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25070 \$153 \$180 \$398 \$179 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25071 \$153 \$180 \$87 \$149 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25073 \$153 \$342 \$57 \$179 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25076 \$153 \$313 \$87 \$178 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25077 \$153 \$229 \$87 \$310 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25078 \$153 \$152 \$23 \$179 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25079 \$16 \$310 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25080 \$16 \$829 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25081 \$16 \$178 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25082 \$153 \$314 \$50 \$309 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25084 \$153 \$230 \$50 \$178 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25085 \$153 \$230 \$549 \$126 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25087 \$153 \$201 \$57 \$126 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25088 \$16 \$276 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25090 \$16 \$310 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25093 \$153 \$261 \$50 \$310 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25095 \$153 \$170 \$23 \$126 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25096 \$153 \$261 \$223 \$126 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25097 \$16 \$149 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25100 \$153 \$262 \$277 \$149 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25102 \$153 \$262 \$398 \$181 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25103 \$153 \$171 \$23 \$181 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25104 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$25105 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$25107 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$25108 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$25109 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$25110 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$25111 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$25113 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$25115 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$25116 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$25117 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$25118 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$25119 \$153 \$7331 \$7319 \$7041 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25121 \$153 \$7355 \$7319 \$6783 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25122 \$153 \$6856 \$7319 \$6981 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25123 \$153 \$7331 \$6996 \$6855 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25125 \$153 \$7393 \$7319 \$6784 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25126 \$16 \$6981 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25127 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$25128 \$153 \$7278 \$7319 \$6907 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25129 \$153 \$7246 \$6794 \$7078 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25130 \$16 \$6784 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25133 \$16 \$6907 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25134 \$153 \$7315 \$7319 \$6792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25136 \$16 \$6915 \$16 \$153 \$7078 VNB sky130_fd_sc_hd__inv_1
X$25137 \$153 \$7280 \$7319 \$6979 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25138 \$153 \$7279 \$6913 \$7078 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25139 \$153 \$7315 \$6719 \$6855 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25140 \$16 \$7378 \$16 \$153 \$6855 VNB sky130_fd_sc_hd__inv_1
X$25142 \$16 \$7381 \$7233 \$7394 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$25143 \$16 \$6979 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25144 \$16 \$7547 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25145 \$153 \$7136 \$7053 \$6784 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25146 \$153 \$7332 \$7053 \$7041 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25147 \$153 \$7332 \$6996 \$7137 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25148 \$16 \$6981 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25149 \$16 \$7041 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25152 \$16 \$7381 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25153 \$16 \$6784 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25154 \$16 \$7333 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25155 \$16 \$7378 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25156 \$16 \$7381 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25157 \$153 \$7395 \$7320 \$7041 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25158 \$16 \$7378 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25159 \$153 \$7334 \$7320 \$6860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25160 \$16 \$7041 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25161 \$16 \$6860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25162 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$25163 \$16 \$6784 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25165 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$25166 \$153 \$6731 \$6732 \$6980 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25167 \$153 \$7282 \$7320 \$6792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25168 \$153 \$7395 \$6996 \$7140 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25169 \$16 \$6783 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25170 \$16 \$6792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25171 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$25172 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$25173 \$153 \$7396 \$7234 \$6981 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25175 \$153 \$7152 \$7234 \$6792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25176 \$153 \$7397 \$7234 \$7041 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25177 \$16 \$6792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25179 \$153 \$7283 \$7234 \$6784 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25182 \$153 \$7398 \$7234 \$6907 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25183 \$153 \$7283 \$6794 \$7141 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25184 \$153 \$7249 \$6995 \$7141 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25186 \$16 \$7071 \$7158 \$7153 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$25187 \$16 \$6907 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25188 \$153 \$7356 \$7235 \$6979 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25189 \$16 \$6784 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25192 \$16 \$6909 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25193 \$16 \$7335 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25194 \$16 \$7154 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25195 \$16 \$7071 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25196 \$153 \$7284 \$7235 \$6783 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25197 \$153 \$7356 \$6995 \$7142 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25198 \$16 \$6979 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25200 \$16 \$6783 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25201 \$153 \$7285 \$7235 \$6784 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25202 \$16 \$7399 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25205 \$153 \$7284 \$6749 \$7142 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25206 \$153 \$7235 \$8365 \$7400 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$25207 \$153 \$7285 \$6794 \$7142 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25208 \$16 \$6981 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25209 \$16 \$6784 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25210 \$16 \$7502 \$16 \$153 \$7142 VNB sky130_fd_sc_hd__inv_1
X$25211 \$16 \$8365 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25213 \$153 \$7401 \$7236 \$6979 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25215 \$153 \$7336 \$7236 \$7041 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25216 \$16 \$6979 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25217 \$153 \$7286 \$7236 \$6860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25218 \$16 \$7041 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25219 \$153 \$7023 \$6913 \$6795 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25221 \$16 \$6784 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25223 \$153 \$7402 \$7337 \$6860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25225 \$153 \$7338 \$7337 \$6784 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25226 \$16 \$6981 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25227 \$16 \$6860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25228 \$16 \$6860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25229 \$16 \$7072 \$7158 \$7287 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$25231 \$153 \$7403 \$7337 \$7041 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25233 \$153 \$7339 \$7337 \$6792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25234 \$16 \$7041 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25236 \$16 \$7379 \$16 \$153 \$7521 VNB sky130_fd_sc_hd__clkbuf_2
X$25237 \$16 \$6792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25238 \$16 \$6784 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25239 \$153 \$153 \$6794 \$7250 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25240 \$153 \$153 \$6732 \$7250 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25242 \$153 \$153 \$6719 \$7250 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25243 \$153 \$153 \$6749 \$7250 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25244 \$16 \$7288 \$16 \$153 \$7250 VNB sky130_fd_sc_hd__clkbuf_2
X$25245 \$153 \$153 \$6913 \$7250 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25246 \$153 \$7073 \$7237 \$7321 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$25247 \$16 \$7545 \$6990 \$7321 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$25248 \$153 \$7370 \$6992 \$7380 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25250 \$153 \$7340 \$7357 \$6862 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25251 \$153 \$7370 \$7357 \$6991 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25252 \$153 \$7221 \$7073 \$6754 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25253 \$16 \$7545 \$16 \$153 \$6982 VNB sky130_fd_sc_hd__inv_1
X$25254 \$16 \$7381 \$16 \$153 \$7380 VNB sky130_fd_sc_hd__inv_1
X$25255 \$16 \$6991 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25257 \$153 \$7191 \$7003 \$6982 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25258 \$16 \$6754 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25259 \$16 \$7381 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25260 \$16 \$6695 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25263 \$153 \$7358 \$7357 \$6771 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25264 \$153 \$7289 \$7073 \$7044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25265 \$153 \$7358 \$6865 \$7380 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25268 \$153 \$7289 \$7006 \$6982 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25269 \$153 \$7404 \$7006 \$7380 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25270 \$16 \$6987 \$6990 \$7160 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$25271 \$16 \$7044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25272 \$16 \$6771 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25273 \$153 \$7341 \$7322 \$6797 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25275 \$153 \$7383 \$6992 \$7382 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25277 \$16 \$6695 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25278 \$153 \$7341 \$6906 \$7382 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25279 \$153 \$7161 \$7322 \$6771 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25280 \$16 \$6797 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25282 \$153 \$7359 \$7322 \$6754 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25283 \$16 \$6771 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25285 \$16 \$6915 \$16 \$153 \$6713 VNB sky130_fd_sc_hd__inv_1
X$25286 \$16 \$7060 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25288 \$153 \$7080 \$7322 \$6862 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25289 \$153 \$7359 \$6756 \$7382 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25290 \$153 \$7405 \$6867 \$7382 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25291 \$16 \$6862 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25292 \$16 \$6989 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25294 \$153 \$7290 \$7323 \$6754 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25295 \$16 \$6754 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25297 \$16 \$8365 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25298 \$16 \$6862 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25300 \$153 \$7406 \$7323 \$6797 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25301 \$16 \$6754 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25303 \$153 \$7005 \$7323 \$7044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25304 \$153 \$7371 \$6324 \$6652 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25305 \$153 \$6870 \$8365 \$7407 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$25307 \$153 \$7223 \$7006 \$6652 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25309 \$16 \$7060 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25310 \$153 \$7360 \$6870 \$7044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25311 \$153 \$7324 \$6870 \$7060 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25314 \$153 \$7324 \$6324 \$6918 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25315 \$153 \$7360 \$7006 \$6918 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25316 \$16 \$7000 \$7163 \$7325 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$25317 \$153 \$7408 \$7006 \$7458 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25318 \$153 \$7238 \$7399 \$7325 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$25320 \$153 \$7409 \$7476 \$6991 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25322 \$16 \$7060 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25323 \$16 \$7044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25324 \$16 \$7156 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25325 \$16 \$6991 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25327 \$153 \$7291 \$7238 \$6754 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25328 \$153 \$7410 \$7238 \$6991 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25329 \$153 \$7291 \$6756 \$7316 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25330 \$16 \$7000 \$16 \$153 \$7316 VNB sky130_fd_sc_hd__inv_1
X$25333 \$16 \$6991 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25334 \$16 \$7000 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25335 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$25336 \$153 \$7292 \$7238 \$6797 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25337 \$153 \$7361 \$7238 \$6771 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25339 \$16 \$6910 \$7163 \$7251 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$25340 \$153 \$7361 \$6865 \$7316 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25343 \$153 \$7292 \$6906 \$7316 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25344 \$16 \$6771 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25346 \$16 \$6935 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25348 \$153 \$7293 \$7252 \$6771 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25349 \$153 \$7362 \$7252 \$7044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25350 \$153 \$7293 \$6865 \$7254 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25351 \$16 \$7044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25353 \$153 \$7362 \$7006 \$7254 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25354 \$16 \$6771 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25356 \$153 \$7363 \$7384 \$6754 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25357 \$16 \$6797 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25358 \$153 \$7166 \$7252 \$7060 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25359 \$153 \$7363 \$6756 \$7411 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25361 \$16 \$6754 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25362 \$16 \$7342 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25363 \$16 \$3418 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25364 \$16 \$3418 \$7342 \$16 \$7412 \$153 VNB sky130_fd_sc_hd__and2_2
X$25366 \$153 \$7294 \$7384 \$7044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25367 \$153 \$7413 \$7384 \$6991 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25368 \$16 \$6991 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25369 \$16 \$6771 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25370 \$153 \$7255 \$6992 \$7254 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25372 \$153 \$7214 \$7003 \$7254 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25373 \$16 \$7060 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25374 \$153 \$7413 \$6992 \$7411 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25376 \$153 \$7295 \$7013 \$7387 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25377 \$16 \$7387 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25378 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$25379 \$153 \$7385 \$7066 \$7296 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25382 \$153 \$7253 \$7013 \$7445 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25383 \$153 \$7364 \$7013 \$7328 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25384 \$16 \$7445 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25386 \$153 \$7343 \$7014 \$7445 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25387 \$16 \$7386 \$16 \$153 \$5932 VNB sky130_fd_sc_hd__inv_1
X$25388 \$16 \$7328 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25389 \$16 \$7445 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25392 \$16 \$7344 \$7633 \$7414 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$25393 \$153 \$7343 \$7327 \$7257 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25394 \$16 \$7344 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25396 \$16 \$7387 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25397 \$153 \$7258 \$7014 \$7387 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25399 \$153 \$7326 \$7014 \$7328 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25401 \$153 \$7326 \$7366 \$7257 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25402 \$16 \$7344 \$16 \$153 \$7257 VNB sky130_fd_sc_hd__inv_1
X$25403 \$16 \$7387 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25404 \$153 \$7259 \$6972 \$7387 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25405 \$153 \$7297 \$6972 \$7328 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25406 \$16 \$7551 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25407 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$25408 \$16 \$7129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25410 \$16 \$7445 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25411 \$153 \$7297 \$7366 \$7146 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25412 \$153 \$7298 \$6972 \$7445 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25414 \$16 \$7350 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25415 \$16 \$7350 \$16 \$153 \$7146 VNB sky130_fd_sc_hd__inv_1
X$25416 \$153 \$7372 \$7066 \$7388 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25417 \$153 \$7298 \$7327 \$7146 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25418 \$153 \$7365 \$7074 \$7387 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25421 \$153 \$7260 \$7482 \$7146 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25423 \$153 \$7261 \$7482 \$7085 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25424 \$153 \$7365 \$7490 \$7085 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25426 \$153 \$7299 \$7074 \$7328 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25427 \$16 \$7328 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25428 \$16 \$7130 \$7633 \$7415 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$25430 \$153 \$7389 \$7065 \$7388 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25431 \$153 \$7299 \$7366 \$7085 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25432 \$16 \$7130 \$16 \$153 \$7085 VNB sky130_fd_sc_hd__inv_1
X$25433 \$16 \$7328 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25434 \$153 \$7416 \$7086 \$7328 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25435 \$16 \$7239 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25436 \$153 \$7300 \$7482 \$6656 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25439 \$153 \$7329 \$7490 \$7112 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25440 \$153 \$7329 \$7086 \$7387 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25442 \$153 \$7301 \$7169 \$7239 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25444 \$153 \$7345 \$7065 \$7317 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25445 \$153 \$7345 \$7169 \$7082 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25447 \$153 \$7367 \$7169 \$7129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25448 \$153 \$7301 \$7482 \$7317 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25450 \$16 \$7445 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25451 \$153 \$7538 \$7170 \$7445 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25452 \$16 \$7082 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25453 \$16 \$7328 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25455 \$153 \$7346 \$7170 \$7328 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25456 \$16 \$7129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25458 \$153 \$7346 \$7366 \$6656 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25460 \$16 \$6656 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25461 \$153 \$7373 \$7066 \$7264 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25462 \$16 \$6656 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25463 \$16 \$7239 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25464 \$153 \$7263 \$7171 \$7239 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25466 \$153 \$7373 \$7171 \$7029 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25467 \$153 \$7262 \$7171 \$7129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25468 \$16 \$7029 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25469 \$16 \$7082 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25470 \$153 \$7374 \$7065 \$7417 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25473 \$153 \$7374 \$7265 \$7082 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25474 \$153 \$7302 \$7265 \$7029 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25476 \$16 \$7387 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25477 \$153 \$7266 \$7366 \$7172 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25478 \$153 \$7047 \$7215 \$7172 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25479 \$153 \$7303 \$7090 \$7387 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25481 \$153 \$7205 \$7065 \$7172 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25482 \$153 \$7304 \$6582 \$7417 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25483 \$153 \$7303 \$7490 \$7172 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25484 \$153 \$7330 \$7090 \$7445 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25485 \$16 \$7445 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25489 \$16 \$7498 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25490 \$153 \$7330 \$7327 \$7172 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25491 \$16 \$7498 \$16 \$153 \$7172 VNB sky130_fd_sc_hd__inv_1
X$25492 \$153 \$7305 \$7482 \$7417 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25493 \$153 \$7216 \$7482 \$7172 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25494 \$16 \$7344 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25495 \$16 \$7344 \$7049 \$7450 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$25496 \$16 \$7386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25497 \$16 \$7347 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25499 \$16 \$7049 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25500 \$16 \$7377 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25501 \$16 \$7484 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25503 \$153 \$7348 \$7173 \$7307 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25504 \$153 \$7418 \$7173 \$7377 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25505 \$153 \$7348 \$7607 \$7093 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25506 \$153 \$7268 \$7180 \$7093 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25508 \$16 \$7307 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25509 \$153 \$7419 \$7173 \$7353 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25512 \$153 \$7269 \$7173 \$7464 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25513 \$153 \$7240 \$8869 \$7349 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$25514 \$16 \$7130 \$7049 \$7349 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$25515 \$16 \$7464 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25517 \$153 \$7175 \$7240 \$7131 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25519 \$153 \$7420 \$7240 \$7307 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25520 \$16 \$7130 \$16 \$153 \$7148 VNB sky130_fd_sc_hd__inv_1
X$25521 \$16 \$7147 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25522 \$16 \$7307 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25524 \$153 \$7421 \$7240 \$7377 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25525 \$153 \$7271 \$7180 \$7148 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25527 \$153 \$7177 \$7241 \$7131 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25528 \$16 \$7131 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25529 \$16 \$7049 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25530 \$16 \$7377 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25531 \$153 \$7422 \$7241 \$7377 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25532 \$153 \$7096 \$7241 \$7174 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25535 \$153 \$7390 \$7639 \$7097 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25537 \$16 \$7350 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25538 \$16 \$7307 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25539 \$16 \$7353 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25541 \$153 \$7368 \$7241 \$7353 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25542 \$153 \$7351 \$7241 \$7307 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25543 \$153 \$7368 \$7375 \$7097 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25545 \$153 \$7273 \$7463 \$7097 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25546 \$16 \$7350 \$16 \$153 \$7097 VNB sky130_fd_sc_hd__inv_1
X$25547 \$16 \$7133 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25549 \$153 \$7423 \$7242 \$7174 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25550 \$153 \$7352 \$7242 \$7133 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25551 \$16 \$5963 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25554 \$16 \$7131 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25555 \$153 \$7352 \$7180 \$7149 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25556 \$16 \$7049 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25557 \$16 \$7131 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25558 \$153 \$7183 \$7243 \$7131 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25559 \$153 \$7423 \$7376 \$7149 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25560 \$153 \$7391 \$7639 \$7392 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25561 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$25562 \$16 \$7174 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25563 \$153 \$7274 \$7463 \$7392 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25566 \$153 \$7354 \$7243 \$7174 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25567 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$25568 \$153 \$7354 \$7376 \$7392 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25569 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$25570 \$16 \$7131 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25571 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$25572 \$153 \$7308 \$7244 \$7131 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25573 \$16 \$7307 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25575 \$153 \$7424 \$7244 \$7307 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25576 \$16 \$7489 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25578 \$16 \$7353 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25580 \$153 \$7425 \$7244 \$7353 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25582 \$153 \$7309 \$7208 \$7217 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25585 \$16 \$7540 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25586 \$16 \$7131 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25587 \$153 \$7310 \$7208 \$7318 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25588 \$16 \$7540 \$7496 \$7426 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$25589 \$16 \$7377 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25590 \$153 \$7427 \$7186 \$7377 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25591 \$153 \$7310 \$7186 \$7131 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25593 \$153 \$7428 \$7186 \$7307 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25594 \$153 \$7311 \$7186 \$7133 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25595 \$153 \$7276 \$7463 \$7318 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25597 \$153 \$5401 \$3142 \$5158 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25598 \$16 \$7614 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25599 \$16 \$7429 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25601 \$16 \$5158 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25602 \$16 \$7353 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25604 \$16 \$7464 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25605 \$16 \$7133 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25606 \$153 \$7430 \$7245 \$7353 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25607 \$153 \$7617 \$7245 \$7133 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25608 \$16 \$7431 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25609 \$16 \$7429 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25611 \$16 \$7377 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25613 \$16 \$7131 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25614 \$16 \$7353 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25615 \$16 \$7133 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25617 \$153 \$7369 \$7245 \$7377 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25618 \$153 \$7309 \$7245 \$7131 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25620 \$153 \$6495 \$5806 \$6924 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25621 \$16 \$6924 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25622 \$153 \$6553 \$5627 \$6924 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25625 \$153 \$7312 \$7187 \$7133 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25627 \$153 \$7432 \$7187 \$7353 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25628 \$153 \$5308 \$3142 \$4963 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25629 \$16 \$4963 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25630 \$153 \$5146 \$4414 \$4963 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25632 \$153 \$7118 \$5806 \$6760 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25635 \$16 \$7464 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25636 \$153 \$7433 \$7187 \$7464 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25637 \$153 \$7313 \$7187 \$7307 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25638 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$25639 \$153 \$6899 \$5635 \$6760 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25640 \$16 \$7307 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25641 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$25643 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$25644 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$25645 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$25646 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$25647 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$25648 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$25649 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$25651 \$153 \$8087 \$8113 \$7041 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25652 \$153 \$8201 \$6930 \$8034 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25653 \$153 \$8087 \$6996 \$8034 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25654 \$153 \$8202 \$6749 \$8034 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25655 \$16 \$6783 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25657 \$153 \$8173 \$8113 \$6907 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25658 \$16 \$6981 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25659 \$16 \$7041 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25661 \$153 \$8033 \$8113 \$6860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25662 \$153 \$8173 \$6913 \$8034 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25663 \$16 \$6860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25664 \$16 \$6907 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25665 \$16 \$6979 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25666 \$153 \$8203 \$6719 \$8034 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25668 \$153 \$8138 \$8113 \$6979 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25669 \$153 \$8138 \$6995 \$8034 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25670 \$16 \$6979 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25671 \$16 \$8167 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25672 \$16 \$8139 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25673 \$153 \$8174 \$8194 \$7816 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25674 \$153 \$7941 \$7784 \$6783 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25676 \$16 \$8139 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25677 \$16 \$8193 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25678 \$153 \$8204 \$6995 \$8206 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25679 \$153 \$8140 \$7784 \$6860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25680 \$16 \$6783 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25681 \$16 \$8114 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25682 \$153 \$8140 \$6732 \$7711 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25683 \$16 \$6860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25684 \$16 \$8114 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25685 \$153 \$8205 \$6930 \$8206 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25687 \$16 \$8003 \$8024 \$8056 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$25688 \$16 \$8423 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25691 \$153 \$8228 \$8115 \$6979 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25692 \$153 \$8035 \$8115 \$6792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25693 \$16 \$6792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25694 \$16 \$6979 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25696 \$16 \$8423 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25697 \$153 \$8141 \$8115 \$6783 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25700 \$153 \$8104 \$8115 \$6981 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25701 \$16 \$6783 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25703 \$153 \$7961 \$6930 \$7587 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25704 \$16 \$6981 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25705 \$16 \$7659 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25706 \$16 \$8144 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25707 \$16 \$7655 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25708 \$153 \$8230 \$8297 \$8229 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$25711 \$16 \$7467 \$16 \$153 \$8024 VNB sky130_fd_sc_hd__clkbuf_2
X$25712 \$153 \$8004 \$7866 \$6784 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25713 \$16 \$8297 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25715 \$16 \$7816 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25716 \$16 \$8144 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25717 \$153 \$8336 \$6732 \$8208 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25718 \$153 \$8104 \$6930 \$8036 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25721 \$153 \$8207 \$8209 \$7816 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25723 \$153 \$7932 \$7866 \$6981 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25724 \$153 \$8175 \$6995 \$8208 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25725 \$153 \$7555 \$6995 \$7608 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25726 \$153 \$8725 \$8737 \$7816 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25728 \$16 \$7973 \$8195 \$8116 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$25730 \$153 \$7866 \$8117 \$8116 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$25731 \$16 \$7973 \$16 \$153 \$7609 VNB sky130_fd_sc_hd__inv_1
X$25732 \$153 \$7701 \$8025 \$8176 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$25733 \$16 \$7816 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25735 \$153 \$8088 \$7701 \$7041 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25736 \$16 \$8118 \$8195 \$8176 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$25737 \$16 \$6979 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25739 \$153 \$7987 \$6749 \$7609 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25740 \$16 \$8118 \$16 \$153 \$7772 VNB sky130_fd_sc_hd__inv_1
X$25741 \$16 \$7041 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25742 \$16 \$7663 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25743 \$16 \$7663 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25744 \$153 \$7966 \$7703 \$6792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25746 \$16 \$6792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25748 \$153 \$7942 \$7703 \$6860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25750 \$16 \$6792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25751 \$16 \$8125 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25752 \$16 \$6860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25753 \$16 \$8061 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25754 \$16 \$6935 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25755 \$153 \$8058 \$6996 \$7768 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25756 \$16 \$8119 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25757 \$16 \$8125 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25758 \$153 \$8210 \$6719 \$8196 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25759 \$153 \$8059 \$6749 \$7768 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25760 \$16 \$8177 \$8195 \$8168 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$25761 \$153 \$7703 \$8061 \$8060 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$25762 \$16 \$7945 \$8169 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$25764 \$153 \$8211 \$6913 \$8196 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25765 \$16 \$8062 \$16 \$153 \$7663 VNB sky130_fd_sc_hd__clkbuf_2
X$25767 \$153 \$8178 \$6995 \$8196 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25768 \$16 \$8063 \$16 \$153 \$8125 VNB sky130_fd_sc_hd__clkbuf_2
X$25769 \$153 \$8120 \$8026 \$8037 \$7989 \$8005 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$25770 \$153 \$7965 \$6794 \$7772 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25772 \$153 \$7988 \$6913 \$7772 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25773 \$153 \$7820 \$6732 \$7772 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25774 \$153 \$7989 \$8005 \$8142 \$8026 \$8037 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$25776 \$16 \$8037 \$8005 \$8026 \$7989 \$16 \$153 \$8233 VNB
+ sky130_fd_sc_hd__and4_2
X$25777 \$16 \$7822 \$16 \$153 \$6915 VNB sky130_fd_sc_hd__clkbuf_2
X$25778 \$153 \$8026 \$8005 \$8143 \$7989 \$8037 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$25779 \$16 \$7888 \$16 \$153 \$7378 VNB sky130_fd_sc_hd__clkbuf_2
X$25780 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25781 \$16 \$8121 \$7226 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$25784 \$16 \$8197 \$16 \$153 \$8001 VNB sky130_fd_sc_hd__clkbuf_2
X$25785 \$16 \$8105 \$16 \$153 \$7922 VNB sky130_fd_sc_hd__clkbuf_2
X$25786 \$153 \$8197 \$8067 \$7990 \$8066 \$8038 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$25787 \$153 \$8105 \$8066 \$7990 \$8038 \$8067 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$25788 \$16 \$7990 \$8067 \$8066 \$8038 \$16 \$153 \$8039 VNB
+ sky130_fd_sc_hd__and4_2
X$25789 \$153 \$8066 \$8067 \$8212 \$8038 \$7990 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$25790 \$16 \$8106 \$16 \$153 \$8144 VNB sky130_fd_sc_hd__clkbuf_2
X$25792 \$153 \$7946 \$7884 \$8145 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$25794 \$16 \$7922 \$7968 \$8068 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$25795 \$16 \$8001 \$7968 \$8145 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$25796 \$16 \$7945 \$6887 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$25797 \$16 \$7945 \$8117 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$25798 \$153 \$8089 \$7946 \$6797 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25799 \$16 \$6862 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25800 \$16 \$8001 \$16 \$153 \$7787 VNB sky130_fd_sc_hd__inv_1
X$25801 \$153 \$8146 \$6992 \$7787 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25803 \$153 \$8213 \$7003 \$8214 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25804 \$153 \$8146 \$7946 \$6991 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25806 \$153 \$8122 \$7946 \$6771 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25807 \$153 \$8089 \$6906 \$7787 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25808 \$16 \$6797 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25809 \$153 \$8069 \$6324 \$7787 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25811 \$153 \$8122 \$6865 \$7787 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25812 \$16 \$6771 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25813 \$16 \$6991 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25814 \$16 \$8114 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25815 \$16 \$7060 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25817 \$153 \$8123 \$8147 \$6754 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25819 \$153 \$8090 \$8147 \$6797 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25821 \$16 \$6754 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25822 \$153 \$8123 \$6756 \$8107 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25823 \$16 \$6797 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25824 \$16 \$7884 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25825 \$16 \$8001 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25826 \$153 \$8179 \$8147 \$6991 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25827 \$153 \$8090 \$6906 \$8107 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25828 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$25830 \$153 \$8179 \$6992 \$8107 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25831 \$16 \$6991 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25834 \$153 \$8305 \$7003 \$8107 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25835 \$153 \$8124 \$7947 \$6862 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25836 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$25837 \$153 \$8124 \$7003 \$8040 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25838 \$16 \$8144 \$7968 \$8235 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$25839 \$153 \$8148 \$7947 \$6754 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25840 \$16 \$6862 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25842 \$16 \$8144 \$16 \$153 \$7718 VNB sky130_fd_sc_hd__inv_1
X$25843 \$16 \$8144 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25845 \$153 \$8148 \$6756 \$8040 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25846 \$16 \$6754 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25847 \$153 \$8149 \$7707 \$6862 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25848 \$16 \$6771 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25850 \$16 \$8169 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25851 \$16 \$7466 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25852 \$153 \$8149 \$7003 \$7718 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25854 \$153 \$8070 \$7006 \$7718 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25855 \$153 \$7684 \$8169 \$8150 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$25856 \$16 \$8177 \$7804 \$8150 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$25857 \$16 \$6862 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25858 \$153 \$8041 \$7684 \$6991 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25859 \$153 \$8215 \$7003 \$8217 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25861 \$153 \$8216 \$6992 \$8217 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25863 \$16 \$7992 \$7804 \$8151 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$25864 \$16 \$6991 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25865 \$153 \$7975 \$7684 \$7060 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25866 \$153 \$7788 \$8119 \$8151 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$25867 \$153 \$8071 \$6867 \$7895 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25868 \$16 \$7060 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25870 \$16 \$7992 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25871 \$16 \$8118 \$7804 \$8091 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$25872 \$153 \$8236 \$6867 \$8218 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25873 \$153 \$8152 \$7788 \$7060 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25874 \$153 \$8338 \$7006 \$8218 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25875 \$16 \$6991 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25876 \$16 \$7060 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25877 \$153 \$8108 \$7788 \$6862 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25878 \$16 \$6862 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25880 \$153 \$8152 \$6324 \$7720 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25881 \$153 \$8339 \$7003 \$8218 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25882 \$153 \$8108 \$7003 \$7720 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25883 \$153 \$8027 \$8061 \$8153 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$25884 \$16 \$8125 \$7804 \$8153 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$25887 \$153 \$8154 \$8027 \$6754 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25888 \$16 \$8061 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25889 \$16 \$8125 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25890 \$16 \$6753 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25892 \$153 \$8154 \$6756 \$7933 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25893 \$153 \$8155 \$8027 \$6916 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25894 \$16 \$6754 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25895 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$25897 \$153 \$8155 \$6867 \$7933 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25898 \$153 \$8042 \$8027 \$6862 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25899 \$16 \$6916 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25900 \$153 \$8180 \$8027 \$6797 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25901 \$16 \$7060 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25902 \$16 \$6862 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25904 \$16 \$7829 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25906 \$153 \$8180 \$6906 \$7933 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25907 \$153 \$8311 \$7006 \$7933 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25908 \$153 \$8170 \$7003 \$8260 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25909 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$25910 \$153 \$153 \$6867 \$7872 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25911 \$16 \$6797 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25912 \$153 \$153 \$7327 \$8219 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25913 \$16 \$16 \$153 VNB sky130_fd_sc_hd__conb_1
X$25914 \$16 \$8126 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25915 \$153 \$153 \$6992 \$7872 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25917 \$153 \$153 \$7366 \$8219 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25918 \$153 \$153 \$7003 \$7872 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25919 \$153 \$153 \$7482 \$8219 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25920 \$153 \$153 \$7066 \$8219 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25921 \$16 \$7003 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25923 \$16 \$8078 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25924 \$153 \$8238 \$8028 \$7445 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25925 \$16 \$7387 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25927 \$153 \$7901 \$8028 \$7129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25928 \$153 \$8072 \$7490 \$7860 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25929 \$16 \$7129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25931 \$153 \$7993 \$7366 \$7860 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25932 \$16 \$7445 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25933 \$16 \$7994 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25934 \$16 \$7029 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25935 \$16 \$7239 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25937 \$153 \$8127 \$7066 \$7860 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25939 \$153 \$8181 \$7874 \$7239 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25940 \$153 \$7832 \$7215 \$7597 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25941 \$153 \$8181 \$7482 \$7924 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25942 \$153 \$8128 \$6582 \$7924 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25943 \$16 \$7386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25946 \$16 \$7387 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25947 \$16 \$8157 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25948 \$153 \$8182 \$7874 \$7387 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25949 \$16 \$7082 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25950 \$153 \$7875 \$7874 \$7082 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25951 \$153 \$8182 \$7490 \$7924 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25952 \$153 \$8129 \$7066 \$7789 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25955 \$153 \$8129 \$7876 \$7029 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25956 \$153 \$7861 \$7876 \$7067 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25957 \$16 \$7029 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25958 \$153 \$8130 \$7065 \$8043 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25959 \$16 \$8220 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25960 \$16 \$7129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25961 \$153 \$8014 \$8183 \$7129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25964 \$153 \$8074 \$7490 \$7789 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25965 \$153 \$8092 \$7876 \$7328 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25966 \$16 \$7328 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25968 \$16 \$8250 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25969 \$153 \$8221 \$6582 \$8043 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25970 \$16 \$8044 \$16 \$153 \$7789 VNB sky130_fd_sc_hd__inv_1
X$25971 \$153 \$8092 \$7366 \$7789 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25974 \$16 \$8136 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25975 \$16 \$7082 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25976 \$153 \$7635 \$8136 \$8240 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$25978 \$16 \$7328 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25979 \$153 \$8045 \$7635 \$7328 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25981 \$16 \$7029 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25982 \$153 \$8223 \$7065 \$8222 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25983 \$16 \$7904 \$16 \$153 \$7571 VNB sky130_fd_sc_hd__inv_1
X$25985 \$16 \$7387 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25986 \$153 \$8158 \$8029 \$7387 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25987 \$153 \$8046 \$8029 \$7029 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25988 \$153 \$8158 \$7490 \$8222 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25990 \$16 \$7445 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25991 \$153 \$8159 \$8029 \$7445 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25994 \$153 \$8159 \$7327 \$8222 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$25995 \$153 \$8015 \$8184 \$7082 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25996 \$153 \$8241 \$8184 \$7129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$25997 \$16 \$7082 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$25998 \$16 \$7129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26002 \$16 \$7239 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26003 \$16 \$7445 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26004 \$153 \$8242 \$8184 \$7445 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26005 \$153 \$8350 \$8184 \$7239 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26006 \$16 \$7915 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26007 \$153 \$7202 \$7215 \$6656 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26008 \$16 \$7067 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26009 \$153 \$8075 \$7327 \$7726 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26012 \$153 \$8243 \$8030 \$7029 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26013 \$153 \$8160 \$8030 \$7067 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26014 \$16 \$7029 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26015 \$153 \$7998 \$7215 \$7726 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26016 \$16 \$7129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26017 \$153 \$8185 \$7215 \$8048 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26019 \$153 \$8161 \$7953 \$7029 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26020 \$153 \$8185 \$7953 \$7129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26021 \$16 \$7082 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26022 \$153 \$8161 \$7066 \$8048 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26023 \$16 \$7076 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26024 \$16 \$7387 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26025 \$153 \$8162 \$7953 \$7387 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26026 \$16 \$7445 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26028 \$153 \$8244 \$8030 \$7445 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26029 \$153 \$8162 \$7490 \$8048 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26031 \$153 \$8132 \$7953 \$7239 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26032 \$153 \$8131 \$7482 \$8264 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26034 \$153 \$8132 \$7482 \$8048 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26036 \$16 \$8163 \$16 \$153 \$7691 VNB sky130_fd_sc_hd__clkbuf_2
X$26037 \$16 \$7559 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26038 \$16 \$8077 \$16 \$153 \$7952 VNB sky130_fd_sc_hd__clkbuf_2
X$26039 \$16 \$7559 \$16 \$153 \$8049 VNB sky130_fd_sc_hd__clkbuf_2
X$26041 \$16 \$6667 \$16 \$153 \$8051 VNB sky130_fd_sc_hd__clkbuf_2
X$26042 \$153 \$7791 \$7792 \$8163 \$7881 \$7880 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$26043 \$16 \$8109 \$8111 \$8110 \$153 \$16 \$8224 VNB sky130_fd_sc_hd__and3_4
X$26044 \$16 \$8109 \$8110 \$8111 \$153 \$8133 \$16 VNB sky130_fd_sc_hd__and3b_4
X$26046 \$16 \$6667 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26048 \$153 \$8111 \$8109 \$8289 \$8110 \$16 \$16 VNB sky130_fd_sc_hd__nor3b_4
X$26049 \$16 \$8078 \$16 \$153 \$8110 VNB sky130_fd_sc_hd__clkbuf_2
X$26051 \$16 \$8050 \$16 \$153 \$7954 VNB sky130_fd_sc_hd__clkbuf_2
X$26052 \$16 \$8134 \$16 \$153 \$7927 VNB sky130_fd_sc_hd__clkbuf_2
X$26054 \$153 \$7048 \$7208 \$7033 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26055 \$16 \$8049 \$16 \$153 \$8225 VNB sky130_fd_sc_hd__clkbuf_2
X$26056 \$16 \$8078 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26057 \$16 \$8078 \$16 \$153 \$8186 VNB sky130_fd_sc_hd__clkbuf_2
X$26060 \$16 \$8112 \$16 \$153 \$8044 VNB sky130_fd_sc_hd__clkbuf_2
X$26061 \$153 \$8198 \$7208 \$7076 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26062 \$153 \$7955 \$7954 \$8079 \$7936 \$7927 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$26063 \$153 \$153 \$7607 \$8186 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26064 \$153 \$153 \$7208 \$8186 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26065 \$153 \$153 \$7180 \$8186 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26066 \$153 \$153 \$7376 \$8186 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26068 \$153 \$153 \$7463 \$8186 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26069 \$16 \$8052 \$16 \$153 \$7667 VNB sky130_fd_sc_hd__clkbuf_2
X$26070 \$16 \$8079 \$16 \$153 \$7709 VNB sky130_fd_sc_hd__clkbuf_2
X$26071 \$153 \$153 \$7639 \$8186 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26072 \$153 \$7938 \$8018 \$7131 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26073 \$16 \$8187 \$8199 \$8247 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$26074 \$16 \$7147 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26075 \$153 \$8188 \$8018 \$7133 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26077 \$16 \$7999 \$16 \$153 \$7386 VNB sky130_fd_sc_hd__clkbuf_2
X$26079 \$153 \$8080 \$7639 \$7928 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26080 \$153 \$8188 \$7180 \$7928 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26081 \$153 \$8094 \$8018 \$7353 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26082 \$16 \$7894 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26083 \$16 \$7894 \$16 \$153 \$7615 VNB sky130_fd_sc_hd__clkbuf_2
X$26085 \$153 \$8226 \$7376 \$7928 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26086 \$153 \$8094 \$7375 \$7928 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26087 \$16 \$8220 \$8199 \$8248 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$26088 \$153 \$7957 \$7862 \$7307 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26090 \$153 \$8249 \$7862 \$7377 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26093 \$16 \$7133 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26094 \$16 \$7904 \$8199 \$8095 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$26095 \$16 \$7147 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26096 \$153 \$8227 \$7463 \$7939 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26097 \$153 \$8096 \$7862 \$7133 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26098 \$153 \$8189 \$8250 \$8251 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$26100 \$153 \$7710 \$8136 \$8095 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$26102 \$153 \$8096 \$7180 \$7939 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26104 \$16 \$7174 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26105 \$153 \$8190 \$8189 \$7174 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26106 \$153 \$8097 \$8189 \$7377 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26107 \$153 \$8190 \$7376 \$8098 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26109 \$153 \$8097 \$7462 \$8098 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26110 \$153 \$8191 \$7607 \$8098 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26111 \$153 \$8082 \$7208 \$8098 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26112 \$16 \$8044 \$16 \$153 \$8098 VNB sky130_fd_sc_hd__inv_1
X$26113 \$153 \$8164 \$8189 \$7147 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26114 \$153 \$7424 \$7607 \$6985 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26116 \$16 \$8044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26118 \$153 \$8164 \$7463 \$8098 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26119 \$153 \$8054 \$8189 \$7133 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26120 \$16 \$7133 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26121 \$153 \$8053 \$8031 \$7133 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26122 \$16 \$7133 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26123 \$16 \$7377 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26124 \$16 \$8266 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26126 \$16 \$8165 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26127 \$16 \$7131 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26128 \$16 \$6985 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26129 \$16 \$7174 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26130 \$16 \$7147 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26131 \$153 \$8813 \$8031 \$7174 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26132 \$153 \$8099 \$8031 \$7147 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26133 \$16 \$7691 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26134 \$16 \$8266 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26135 \$16 \$8135 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26137 \$16 \$7131 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26138 \$16 \$7133 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26139 \$16 \$7147 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26141 \$153 \$8166 \$8200 \$7147 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26143 \$153 \$8171 \$8200 \$7133 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26144 \$16 \$7174 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26145 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$26146 \$153 \$7700 \$7639 \$7882 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26147 \$16 \$7131 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26148 \$153 \$8172 \$8200 \$7131 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26150 \$153 \$8100 \$8200 \$7174 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26151 \$153 \$7699 \$7376 \$7882 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26152 \$16 \$8359 \$8032 \$8137 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$26153 \$153 \$7430 \$7375 \$7217 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26154 \$16 \$7133 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26155 \$153 \$8081 \$7863 \$7133 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26157 \$16 \$7464 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26159 \$16 \$8473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26160 \$153 \$7515 \$7607 \$7217 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26161 \$16 \$8101 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26162 \$16 \$8359 \$16 \$153 \$7076 VNB sky130_fd_sc_hd__inv_1
X$26163 \$153 \$7232 \$7376 \$7217 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26164 \$16 \$8359 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26166 \$153 \$7917 \$7375 \$7782 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26167 \$16 \$8265 \$8032 \$8253 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$26169 \$16 \$8032 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26172 \$16 \$7133 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26173 \$16 \$7147 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26174 \$153 \$8192 \$7960 \$7133 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26175 \$153 \$8102 \$7960 \$7147 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26176 \$16 \$8265 \$16 \$153 \$7033 VNB sky130_fd_sc_hd__inv_1
X$26177 \$153 \$7842 \$7180 \$7782 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26178 \$16 \$8265 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26179 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$26181 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$26182 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$26183 \$16 \$7174 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26184 \$16 \$7464 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26185 \$153 \$8103 \$7960 \$7464 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26186 \$16 \$7307 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26187 \$153 \$8254 \$7960 \$7307 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26188 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$26189 \$153 \$7583 \$7180 \$7763 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26192 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$26194 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$26195 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$26196 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$26197 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$26198 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$26200 \$153 \$1976 \$2193 \$1687 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26201 \$153 \$1684 \$2193 \$1980 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26202 \$16 \$1687 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26203 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$26204 \$16 \$1980 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26205 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$26207 \$153 \$2209 \$1792 \$2110 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26210 \$153 \$2286 \$1943 \$2110 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26211 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$26212 \$153 \$2134 \$1873 \$2024 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26213 \$153 \$2287 \$1547 \$2110 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26214 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$26215 \$153 \$2969 \$2064 \$2110 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26216 \$16 \$2024 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26219 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$26220 \$16 \$2180 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26221 \$16 \$710 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26222 \$153 \$2248 \$1774 \$1942 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26223 \$153 \$2213 \$1774 \$2024 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26224 \$16 \$2180 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26226 \$153 \$1788 \$1774 \$2180 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26227 \$16 \$1942 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26228 \$16 \$1430 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26231 \$16 \$585 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26233 \$16 \$1596 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26234 \$153 \$2212 \$1763 \$2024 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26235 \$153 \$2415 \$1547 \$2179 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26236 \$16 \$2180 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26237 \$16 \$2024 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26238 \$153 \$2274 \$2210 \$1669 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26239 \$16 \$582 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26240 \$16 \$754 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26242 \$153 \$2136 \$1763 \$1795 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26243 \$153 \$2322 \$2064 \$1669 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26244 \$153 \$2324 \$1547 \$1669 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26245 \$153 \$2211 \$1943 \$1789 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26246 \$16 \$1795 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26247 \$16 \$1522 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26248 \$16 \$1687 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26249 \$153 \$2212 \$2210 \$1789 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26250 \$16 \$2006 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26252 \$153 \$2288 \$1888 \$2006 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26253 \$153 \$2136 \$1815 \$1789 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26254 \$153 \$2213 \$2210 \$1537 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26255 \$153 \$2248 \$2064 \$1537 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26256 \$16 \$430 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26257 \$153 \$2288 \$1943 \$1861 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26258 \$16 \$280 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26260 \$153 \$2097 \$1963 \$2180 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26262 \$153 \$2138 \$2210 \$1793 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26263 \$153 \$2249 \$1815 \$2275 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26264 \$153 \$2035 \$1963 \$1942 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26265 \$16 \$2180 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26268 \$153 \$2066 \$2009 \$1793 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26269 \$16 \$1942 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26271 \$153 \$2214 \$1766 \$2024 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26272 \$153 \$2250 \$2064 \$2181 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26273 \$16 \$1430 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26274 \$16 \$1430 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26276 \$16 \$280 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26277 \$16 \$2180 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26278 \$153 \$2214 \$2210 \$1767 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26279 \$16 \$2024 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26281 \$153 \$2087 \$2252 \$1767 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26282 \$153 \$2354 \$1659 \$2215 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$26283 \$16 \$899 \$1522 \$2215 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$26284 \$16 \$899 \$16 \$153 \$2181 VNB sky130_fd_sc_hd__inv_1
X$26285 \$153 \$2141 \$1675 \$2180 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26286 \$153 \$2289 \$2009 \$2181 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26289 \$16 \$1658 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26290 \$153 \$2140 \$2064 \$1796 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26291 \$153 \$2067 \$1943 \$1796 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26292 \$153 \$2290 \$1047 \$2251 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$26293 \$153 \$2141 \$2252 \$1796 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26294 \$16 \$2180 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26295 \$16 \$2024 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26296 \$16 \$849 \$1430 \$2251 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$26299 \$153 \$2216 \$1676 \$2180 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26300 \$16 \$1687 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26301 \$153 \$2243 \$1815 \$2219 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26302 \$153 \$2216 \$2252 \$1670 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26303 \$16 \$2180 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26304 \$16 \$2024 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26306 \$153 \$2243 \$2194 \$1795 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26307 \$16 \$1430 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26308 \$16 \$1047 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26312 \$153 \$2291 \$2210 \$2219 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26314 \$16 \$1687 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26315 \$153 \$2292 \$2194 \$2180 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26316 \$153 \$2217 \$2194 \$1687 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26317 \$153 \$2293 \$2194 \$2006 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26319 \$153 \$2143 \$2064 \$1671 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26321 \$16 \$652 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26322 \$16 \$652 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26323 \$153 \$2194 \$685 \$2218 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$26324 \$153 \$2068 \$2009 \$1671 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26325 \$16 \$652 \$2647 \$2218 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$26327 \$16 \$2182 \$16 \$153 \$691 VNB sky130_fd_sc_hd__clkbuf_2
X$26328 \$153 \$2253 \$2194 \$1658 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26329 \$16 \$2145 \$16 \$153 \$585 VNB sky130_fd_sc_hd__clkbuf_2
X$26330 \$16 \$652 \$16 \$153 \$2219 VNB sky130_fd_sc_hd__inv_1
X$26331 \$16 \$2069 \$16 \$153 \$849 VNB sky130_fd_sc_hd__clkbuf_2
X$26333 \$16 \$2195 \$16 \$153 \$2420 VNB sky130_fd_sc_hd__clkbuf_2
X$26334 \$153 \$2253 \$1547 \$2219 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26335 \$16 \$2195 \$16 \$153 \$2038 VNB sky130_fd_sc_hd__clkbuf_2
X$26336 \$16 \$2113 \$16 \$153 \$1875 VNB sky130_fd_sc_hd__clkbuf_2
X$26337 \$16 \$1980 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26340 \$153 \$2220 \$2183 \$2294 \$2196 \$16 \$16 VNB sky130_fd_sc_hd__nor3b_4
X$26341 \$16 \$2183 \$2196 \$2220 \$153 \$2197 \$16 VNB sky130_fd_sc_hd__and3b_4
X$26342 \$16 \$531 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26343 \$153 \$1875 \$2038 \$2115 \$1863 \$1842 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$26344 \$16 \$1354 \$16 \$153 \$2196 VNB sky130_fd_sc_hd__clkbuf_2
X$26345 \$16 \$2276 \$16 \$153 \$2435 VNB sky130_fd_sc_hd__clkbuf_2
X$26346 \$16 \$2197 \$16 \$153 \$1842 VNB sky130_fd_sc_hd__clkbuf_2
X$26347 \$16 \$585 \$1292 \$2295 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$26348 \$16 \$2070 \$16 \$153 \$1291 VNB sky130_fd_sc_hd__clkbuf_2
X$26350 \$16 \$1037 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26351 \$153 \$2221 \$2039 \$2199 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26352 \$153 \$2146 \$2039 \$1965 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26353 \$16 \$2296 \$16 \$153 \$652 VNB sky130_fd_sc_hd__clkbuf_2
X$26354 \$153 \$2146 \$1806 \$1944 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26355 \$153 \$2297 \$2039 \$2089 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26357 \$153 \$2221 \$2184 \$1944 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26358 \$153 \$2254 \$2039 \$2042 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26359 \$153 \$2088 \$2184 \$1864 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26361 \$153 \$2147 \$2039 \$2043 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26362 \$16 \$2089 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26363 \$16 \$2042 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26365 \$153 \$2254 \$1924 \$1944 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26366 \$153 \$2147 \$1954 \$1944 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26367 \$16 \$2043 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26368 \$16 \$2042 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26369 \$16 \$1805 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26370 \$16 \$2634 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26371 \$153 \$2072 \$1954 \$1864 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26372 \$153 \$2298 \$2244 \$1805 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26373 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$26376 \$16 \$430 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26377 \$153 \$2148 \$2026 \$1483 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26378 \$153 \$2198 \$2244 \$1845 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26379 \$153 \$2244 \$430 \$2150 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$26380 \$16 \$582 \$16 \$153 \$2299 VNB sky130_fd_sc_hd__inv_1
X$26381 \$16 \$1965 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26382 \$16 \$1845 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26383 \$153 \$2149 \$2184 \$1483 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26385 \$16 \$582 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26386 \$16 \$582 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26387 \$16 \$279 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26388 \$153 \$2041 \$1921 \$2089 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26389 \$16 \$1923 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26390 \$153 \$2300 \$1921 \$1845 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26391 \$16 \$2089 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26392 \$153 \$2298 \$1703 \$2299 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26393 \$16 \$710 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26396 \$153 \$2198 \$1471 \$2299 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26397 \$16 \$1845 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26398 \$16 \$1966 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26399 \$16 \$279 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26401 \$153 \$2301 \$1697 \$2199 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26402 \$153 \$2118 \$1697 \$2089 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26403 \$16 \$2199 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26404 \$16 \$2089 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26406 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$26407 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$26408 \$16 \$2362 \$16 \$153 \$1292 VNB sky130_fd_sc_hd__clkbuf_2
X$26409 \$153 \$2222 \$1820 \$2089 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26410 \$153 \$2224 \$1820 \$2042 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26411 \$16 \$849 \$1292 \$2223 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$26412 \$153 \$2222 \$2026 \$1844 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26414 \$153 \$2102 \$1820 \$2199 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26415 \$16 \$2042 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26416 \$16 \$1067 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26418 \$16 \$2199 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26419 \$153 \$2255 \$2277 \$2042 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26420 \$153 \$2224 \$1924 \$1844 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26421 \$16 \$849 \$16 \$153 \$2152 VNB sky130_fd_sc_hd__inv_1
X$26423 \$153 \$2153 \$1700 \$2199 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26425 \$153 \$2255 \$1924 \$2152 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26426 \$16 \$2042 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26428 \$153 \$2185 \$2277 \$1965 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26429 \$153 \$2153 \$2184 \$1822 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26430 \$16 \$2199 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26434 \$153 \$2185 \$1806 \$2152 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26435 \$153 \$2256 \$2277 \$1845 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26436 \$16 \$899 \$1966 \$2329 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$26437 \$153 \$2225 \$2200 \$1923 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26438 \$153 \$2256 \$1471 \$2152 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26441 \$16 \$899 \$16 \$153 \$2186 VNB sky130_fd_sc_hd__inv_1
X$26442 \$16 \$1923 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26444 \$16 \$1965 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26445 \$153 \$2074 \$1924 \$1752 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26447 \$153 \$2257 \$2200 \$2089 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26448 \$153 \$2330 \$1806 \$2186 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26449 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$26450 \$153 \$2257 \$2026 \$2186 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26453 \$153 \$2226 \$1780 \$2042 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26454 \$16 \$2089 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26456 \$153 \$1967 \$685 \$2302 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$26457 \$153 \$2226 \$1924 \$1704 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26458 \$16 \$2042 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26459 \$16 \$685 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26460 \$16 \$2089 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26462 \$16 \$2199 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26463 \$16 \$652 \$16 \$153 \$2028 VNB sky130_fd_sc_hd__inv_1
X$26465 \$153 \$2121 \$1967 \$2199 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26466 \$153 \$2227 \$1967 \$2042 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26468 \$16 \$2042 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26469 \$153 \$2227 \$1924 \$2028 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26471 \$16 \$2043 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26472 \$153 \$2258 \$1967 \$2043 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26475 \$153 \$2158 \$1967 \$2089 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26476 \$153 \$2258 \$1954 \$2028 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26477 \$153 \$2158 \$2026 \$2028 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26478 \$153 \$2259 \$1613 \$2278 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26479 \$153 \$2157 \$1471 \$2028 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26481 \$153 \$2259 \$2279 \$1969 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26482 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$26484 \$153 \$2159 \$1876 \$2105 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26486 \$153 \$2246 \$2279 \$1878 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26489 \$153 \$2159 \$2438 \$1540 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26490 \$153 \$2279 \$558 \$2304 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$26491 \$153 \$2246 \$1868 \$2278 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26492 \$153 \$2046 \$1781 \$2104 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26493 \$153 \$2303 \$1558 \$2161 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26495 \$153 \$2332 \$2092 \$2278 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26496 \$16 \$2105 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26497 \$16 \$2098 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26498 \$153 \$2260 \$2103 \$2098 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26499 \$16 \$1878 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26500 \$153 \$2228 \$2103 \$2105 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26501 \$153 \$2305 \$2103 \$2016 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26503 \$153 \$2162 \$1868 \$2078 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26504 \$16 \$2016 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26506 \$153 \$2201 \$2103 \$1879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26507 \$153 \$2228 \$2438 \$2078 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26508 \$16 \$1879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26509 \$16 \$1969 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26510 \$16 \$1756 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26511 \$153 \$2201 \$1558 \$2078 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26513 \$153 \$2306 \$1712 \$2078 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26515 \$153 \$2307 \$2202 \$1756 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26516 \$153 \$2229 \$2202 \$1969 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26517 \$16 \$1969 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26518 \$16 \$2016 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26521 \$16 \$354 \$1968 \$2261 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$26522 \$153 \$2049 \$1900 \$2016 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26523 \$153 \$2202 \$674 \$2261 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$26524 \$153 \$1615 \$389 \$1811 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26525 \$153 \$2229 \$1613 \$2280 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26526 \$16 \$2105 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26527 \$153 \$2050 \$1880 \$2105 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26529 \$153 \$2308 \$1558 \$2280 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26530 \$16 \$354 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26532 \$16 \$1969 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26533 \$153 \$2163 \$2092 \$1674 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26534 \$153 \$2262 \$2309 \$1969 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26535 \$16 \$1518 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26536 \$16 \$1929 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26538 \$16 \$798 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26540 \$153 \$2164 \$1993 \$1674 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26541 \$153 \$2309 \$948 \$2165 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$26542 \$16 \$2104 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26543 \$153 \$2123 \$1928 \$2104 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26544 \$153 \$2262 \$1613 \$2334 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26545 \$16 \$1878 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26547 \$16 \$948 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26548 \$153 \$2263 \$2310 \$1878 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26549 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$26550 \$16 \$2016 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26551 \$153 \$1714 \$1928 \$2016 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26553 \$153 \$2310 \$116 \$2311 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$26555 \$16 \$116 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26557 \$153 \$2230 \$1712 \$2187 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26558 \$153 \$2312 \$2310 \$1969 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26559 \$16 \$1969 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26560 \$16 \$2104 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26561 \$153 \$2203 \$1903 \$2104 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26562 \$153 \$2081 \$1715 \$1759 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26565 \$16 \$2016 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26566 \$153 \$2203 \$2092 \$1759 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26567 \$16 \$80 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26569 \$16 \$1969 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26570 \$153 \$2231 \$2368 \$1969 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26572 \$16 \$1456 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26573 \$16 \$1456 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26574 \$16 \$2104 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26576 \$153 \$2247 \$1993 \$1996 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26577 \$153 \$2247 \$1854 \$2098 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26579 \$153 \$2231 \$1613 \$2188 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26580 \$153 \$2167 \$1854 \$2016 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26581 \$16 \$2098 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26582 \$16 \$2016 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26584 \$16 \$724 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26585 \$153 \$2281 \$1868 \$2188 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26586 \$153 \$2167 \$1715 \$1996 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26589 \$153 \$1854 \$895 \$2313 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$26590 \$16 \$2168 \$16 \$153 \$2232 VNB sky130_fd_sc_hd__clkbuf_2
X$26591 \$153 \$2054 \$1831 \$1812 \$1782 \$1970 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$26593 \$16 \$2189 \$16 \$153 \$1831 VNB sky130_fd_sc_hd__clkbuf_2
X$26594 \$16 \$2204 \$16 \$153 \$1970 VNB sky130_fd_sc_hd__clkbuf_2
X$26595 \$16 \$1812 \$1831 \$1782 \$1970 \$16 \$153 \$2124 VNB
+ sky130_fd_sc_hd__and4_2
X$26597 \$16 \$2349 \$2315 \$2370 \$153 \$16 \$2314 VNB sky130_fd_sc_hd__and3_4
X$26599 \$16 \$2233 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26600 \$16 \$2204 \$16 \$153 \$1905 VNB sky130_fd_sc_hd__clkbuf_2
X$26601 \$16 \$2233 \$16 \$153 \$2315 VNB sky130_fd_sc_hd__clkbuf_2
X$26602 \$16 \$2126 \$16 \$153 \$1883 VNB sky130_fd_sc_hd__clkbuf_2
X$26603 \$16 \$2463 \$16 \$153 \$1855 VNB sky130_fd_sc_hd__clkbuf_2
X$26604 \$16 \$2189 \$16 \$153 \$1971 VNB sky130_fd_sc_hd__clkbuf_2
X$26606 \$153 \$2316 \$558 \$2264 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$26607 \$153 \$1883 \$1971 \$2205 \$1905 \$1855 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$26608 \$16 \$1855 \$1971 \$1883 \$1905 \$16 \$153 \$2127 VNB
+ sky130_fd_sc_hd__and4_2
X$26610 \$16 \$594 \$1972 \$2264 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$26611 \$16 \$2205 \$16 \$153 \$354 VNB sky130_fd_sc_hd__clkbuf_2
X$26613 \$153 \$2128 \$1906 \$2085 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26614 \$153 \$2234 \$1906 \$2191 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26615 \$16 \$2191 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26616 \$153 \$2234 \$2267 \$1999 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26617 \$16 \$2085 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26620 \$153 \$2235 \$1906 \$2093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26621 \$16 \$2191 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26622 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$26623 \$16 \$1585 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26624 \$153 \$2235 \$2265 \$1999 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26625 \$16 \$2093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26626 \$16 \$2093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26627 \$153 \$2338 \$2265 \$2402 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26629 \$16 \$2085 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26630 \$153 \$2190 \$1974 \$2192 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26632 \$153 \$2317 \$1974 \$2085 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26633 \$153 \$2190 \$2269 \$2129 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26635 \$16 \$2191 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26636 \$153 \$2266 \$1974 \$2191 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26637 \$16 \$2192 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26639 \$16 \$2031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26641 \$16 \$2093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26643 \$153 \$2236 \$1974 \$2093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26644 \$153 \$2266 \$2267 \$2129 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26645 \$16 \$354 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26646 \$153 \$2236 \$2265 \$2129 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26647 \$16 \$2031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26648 \$153 \$2237 \$1909 \$2031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26650 \$16 \$674 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26653 \$16 \$2085 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26654 \$153 \$2318 \$1909 \$2085 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26655 \$153 \$2058 \$674 \$2108 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$26656 \$16 \$798 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26657 \$16 \$856 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26659 \$153 \$2171 \$2265 \$2172 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26660 \$16 \$798 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26661 \$16 \$2191 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26663 \$153 \$2238 \$2058 \$2191 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26664 \$153 \$2268 \$2099 \$2031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26665 \$16 \$798 \$16 \$153 \$2239 VNB sky130_fd_sc_hd__inv_1
X$26666 \$153 \$2268 \$1936 \$2239 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26667 \$153 \$2240 \$2058 \$2192 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26669 \$153 \$2238 \$2267 \$2172 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26670 \$16 \$2192 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26671 \$153 \$2173 \$2099 \$1860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26672 \$153 \$2240 \$2269 \$2172 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26674 \$153 \$2341 \$2269 \$2239 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26675 \$16 \$829 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26678 \$16 \$2192 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26679 \$153 \$2173 \$2000 \$2239 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26680 \$153 \$2270 \$1886 \$2192 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26682 \$153 \$2175 \$1886 \$2093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26683 \$153 \$2270 \$2269 \$2020 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26684 \$153 \$2175 \$2265 \$2020 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26687 \$153 \$2206 \$1886 \$2191 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26688 \$16 \$2191 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26689 \$16 \$151 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26691 \$16 \$80 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26692 \$153 \$2206 \$2267 \$2020 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26693 \$153 \$2632 \$2271 \$2282 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26695 \$16 \$2093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26696 \$153 \$2319 \$2271 \$2020 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26697 \$16 \$2192 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26699 \$153 \$2060 \$2004 \$2192 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26700 \$153 \$2283 \$2086 \$2282 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26701 \$16 \$1600 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26702 \$16 \$2191 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26703 \$16 \$723 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26704 \$153 \$2241 \$2004 \$2191 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26705 \$153 \$2272 \$2271 \$1872 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26707 \$16 \$2085 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26709 \$153 \$2241 \$2267 \$1940 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26710 \$153 \$2176 \$2004 \$2085 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26711 \$16 \$2085 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26712 \$16 \$276 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26713 \$153 \$2320 \$2271 \$2284 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26714 \$16 \$2191 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26715 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$26716 \$153 \$2177 \$2265 \$1872 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26718 \$153 \$2176 \$2271 \$1940 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26719 \$16 \$1860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26720 \$16 \$1973 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26722 \$153 \$2496 \$2000 \$2032 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26723 \$16 \$2031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26724 \$153 \$1916 \$1938 \$2031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26725 \$153 \$2285 \$2056 \$2284 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26728 \$153 \$2242 \$2056 \$2178 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26729 \$16 \$1960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26730 \$153 \$2273 \$2376 \$1960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26731 \$153 \$2207 \$2086 \$2032 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26732 \$153 \$2208 \$1936 \$2284 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26733 \$153 \$2321 \$2269 \$2284 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26735 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$26736 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$26738 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$26739 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$26740 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$26741 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$26742 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$26743 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$26745 \$153 \$529 \$511 \$504 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26746 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$26748 \$153 \$529 \$561 \$598 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26750 \$16 \$504 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26752 \$16 \$17 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26753 \$153 \$617 \$511 \$58 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26754 \$153 \$530 \$511 \$395 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26755 \$153 \$315 \$394 \$88 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26756 \$16 \$395 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26757 \$16 \$264 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26758 \$16 \$531 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26759 \$16 \$503 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26760 \$16 \$58 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26762 \$16 \$264 \$503 \$448 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$26763 \$153 \$618 \$511 \$184 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26765 \$153 \$449 \$377 \$598 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26766 \$153 \$532 \$65 \$504 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26767 \$16 \$184 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26769 \$153 \$532 \$561 \$89 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26771 \$153 \$65 \$1596 \$450 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$26772 \$16 \$504 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26773 \$153 \$429 \$65 \$395 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26774 \$16 \$1596 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26776 \$153 \$562 \$661 \$249 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26777 \$16 \$395 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26778 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$26781 \$153 \$452 \$182 \$419 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26782 \$153 \$562 \$377 \$649 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26783 \$153 \$451 \$561 \$94 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26784 \$153 \$452 \$349 \$94 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26785 \$16 \$754 \$503 \$599 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$26787 \$16 \$279 \$537 \$533 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$26789 \$153 \$182 \$430 \$619 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$26790 \$153 \$500 \$234 \$96 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26791 \$153 \$500 \$66 \$263 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26792 \$16 \$582 \$16 \$153 \$94 VNB sky130_fd_sc_hd__inv_1
X$26794 \$153 \$620 \$66 \$504 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26796 \$16 \$263 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26797 \$16 \$504 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26798 \$153 \$206 \$59 \$96 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26799 \$153 \$554 \$66 \$395 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26800 \$16 \$279 \$16 \$153 \$96 VNB sky130_fd_sc_hd__inv_1
X$26802 \$16 \$503 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26803 \$153 \$455 \$67 \$504 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26804 \$16 \$280 \$503 \$621 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$26807 \$153 \$512 \$67 \$419 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26809 \$153 \$512 \$349 \$270 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26810 \$153 \$455 \$561 \$270 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26811 \$16 \$323 \$503 \$622 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$26812 \$16 \$280 \$16 \$153 \$270 VNB sky130_fd_sc_hd__inv_1
X$26813 \$153 \$563 \$68 \$504 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26814 \$16 \$504 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26816 \$153 \$534 \$68 \$419 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26817 \$153 \$563 \$561 \$98 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26818 \$153 \$534 \$349 \$98 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26819 \$16 \$323 \$16 \$153 \$98 VNB sky130_fd_sc_hd__inv_1
X$26820 \$16 \$504 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26821 \$16 \$419 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26822 \$16 \$323 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26825 \$153 \$513 \$190 \$504 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26827 \$16 \$503 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26828 \$153 \$564 \$349 \$765 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26829 \$16 \$17 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26830 \$16 \$356 \$503 \$565 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$26831 \$16 \$504 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26832 \$153 \$456 \$349 \$100 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26833 \$153 \$69 \$535 \$565 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$26836 \$153 \$513 \$561 \$100 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26837 \$16 \$380 \$537 \$623 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$26838 \$16 \$535 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26840 \$153 \$566 \$69 \$504 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26841 \$16 \$380 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26842 \$153 \$458 \$69 \$419 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26845 \$153 \$566 \$561 \$101 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26846 \$16 \$419 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26847 \$153 \$536 \$583 \$419 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26849 \$153 \$624 \$583 \$249 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26850 \$153 \$457 \$394 \$101 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26851 \$16 \$351 \$537 \$514 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$26853 \$153 \$70 \$505 \$514 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$26855 \$153 \$625 \$583 \$58 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26856 \$16 \$537 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26858 \$16 \$263 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26859 \$153 \$459 \$394 \$172 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26860 \$16 \$58 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26861 \$16 \$505 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26862 \$16 \$351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26863 \$16 \$249 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26864 \$153 \$431 \$506 \$263 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26866 \$153 \$515 \$506 \$249 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26867 \$16 \$351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26868 \$16 \$715 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26870 \$153 \$515 \$377 \$432 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26871 \$16 \$1173 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26872 \$16 \$584 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26873 \$16 \$58 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26874 \$153 \$567 \$506 \$58 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26876 \$16 \$716 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26877 \$16 \$1596 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26878 \$16 \$531 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26879 \$153 \$516 \$59 \$432 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26880 \$153 \$567 \$30 \$432 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26881 \$153 \$420 \$1596 \$517 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$26882 \$16 \$585 \$555 \$517 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$26883 \$16 \$555 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26885 \$153 \$538 \$420 \$293 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26886 \$153 \$626 \$586 \$293 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26887 \$153 \$461 \$346 \$271 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26888 \$16 \$293 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26889 \$16 \$585 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26890 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$26891 \$153 \$568 \$586 \$73 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26892 \$16 \$293 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26894 \$153 \$538 \$35 \$271 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26895 \$153 \$462 \$253 \$271 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26896 \$153 \$568 \$215 \$641 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26897 \$153 \$434 \$420 \$60 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26898 \$16 \$73 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26900 \$16 \$754 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26901 \$16 \$662 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26904 \$16 \$555 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26905 \$16 \$754 \$555 \$569 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$26906 \$153 \$463 \$347 \$271 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26907 \$153 \$74 \$662 \$569 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$26908 \$153 \$518 \$347 \$641 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26909 \$153 \$570 \$74 \$358 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26910 \$16 \$430 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26911 \$16 \$754 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26913 \$153 \$539 \$74 \$212 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26914 \$153 \$464 \$346 \$175 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26915 \$153 \$540 \$185 \$187 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26916 \$153 \$539 \$347 \$175 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26919 \$153 \$192 \$541 \$466 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$26920 \$153 \$465 \$54 \$175 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26921 \$153 \$467 \$347 \$105 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26922 \$16 \$358 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26923 \$153 \$571 \$587 \$293 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26924 \$16 \$187 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26925 \$16 \$541 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26926 \$16 \$279 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26928 \$16 \$279 \$16 \$153 \$186 VNB sky130_fd_sc_hd__inv_1
X$26929 \$153 \$542 \$192 \$209 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26930 \$153 \$571 \$35 \$600 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26931 \$153 \$24 \$1525 \$468 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$26932 \$153 \$519 \$253 \$105 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26935 \$153 \$469 \$24 \$293 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26936 \$16 \$1525 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26938 \$153 \$572 \$587 \$212 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26939 \$153 \$469 \$35 \$325 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26940 \$16 \$212 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26941 \$153 \$53 \$535 \$601 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$26942 \$16 \$187 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26944 \$153 \$470 \$54 \$325 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26945 \$153 \$471 \$253 \$325 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26946 \$16 \$293 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26947 \$153 \$472 \$53 \$209 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26948 \$153 \$542 \$346 \$186 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26949 \$16 \$356 \$16 \$153 \$176 VNB sky130_fd_sc_hd__inv_1
X$26951 \$153 \$472 \$346 \$176 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26953 \$153 \$383 \$54 \$176 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26954 \$16 \$209 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26955 \$16 \$356 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26957 \$16 \$684 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26958 \$153 \$193 \$684 \$543 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$26959 \$16 \$380 \$507 \$543 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$26960 \$16 \$358 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26961 \$16 \$380 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26964 \$16 \$507 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26966 \$16 \$351 \$507 \$520 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$26967 \$16 \$380 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26968 \$153 \$194 \$505 \$520 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$26969 \$16 \$507 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26971 \$153 \$627 \$521 \$212 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26972 \$153 \$384 \$346 \$20 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26973 \$16 \$212 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26975 \$16 \$505 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26976 \$16 \$1332 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26977 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$26979 \$153 \$628 \$521 \$60 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26980 \$153 \$544 \$521 \$18 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26981 \$153 \$214 \$346 \$188 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26982 \$16 \$60 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26983 \$16 \$18 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26984 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$26986 \$153 \$385 \$347 \$188 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26987 \$153 \$628 \$104 \$769 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26988 \$153 \$473 \$35 \$188 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26989 \$16 \$293 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26990 \$153 \$629 \$421 \$293 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26992 \$153 \$435 \$421 \$60 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$26994 \$153 \$522 \$215 \$436 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26995 \$16 \$588 \$16 \$153 \$436 VNB sky130_fd_sc_hd__inv_1
X$26996 \$16 \$73 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26997 \$16 \$209 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$26998 \$153 \$474 \$54 \$436 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$26999 \$153 \$573 \$421 \$209 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27000 \$16 \$588 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27004 \$153 \$475 \$347 \$436 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27005 \$153 \$573 \$346 \$436 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27006 \$153 \$386 \$253 \$329 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27007 \$153 \$602 \$253 \$436 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27008 \$153 \$545 \$422 \$241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27009 \$16 \$241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27012 \$153 \$40 \$21 \$352 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27014 \$16 \$145 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27015 \$153 \$630 \$422 \$145 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27017 \$16 \$79 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27019 \$153 \$546 \$422 \$79 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27020 \$153 \$422 \$558 \$574 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$27021 \$153 \$478 \$44 \$501 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27022 \$16 \$594 \$397 \$574 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$27023 \$16 \$79 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27024 \$16 \$241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27027 \$153 \$479 \$407 \$79 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27028 \$153 \$557 \$407 \$241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27029 \$153 \$546 \$112 \$501 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27030 \$153 \$330 \$266 \$111 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27031 \$153 \$141 \$112 \$111 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27033 \$153 \$603 \$389 \$604 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27034 \$153 \$589 \$353 \$604 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27035 \$16 \$397 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27036 \$16 \$438 \$397 \$523 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$27037 \$153 \$77 \$631 \$523 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$27038 \$16 \$399 \$16 \$153 \$604 VNB sky130_fd_sc_hd__inv_1
X$27041 \$16 \$631 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27042 \$16 \$79 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27043 \$153 \$575 \$590 \$79 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27045 \$16 \$424 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27046 \$153 \$480 \$77 \$424 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27047 \$153 \$575 \$112 \$605 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27050 \$16 \$438 \$16 \$153 \$113 VNB sky130_fd_sc_hd__inv_1
X$27051 \$153 \$480 \$353 \$113 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27053 \$153 \$78 \$674 \$548 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$27054 \$16 \$354 \$397 \$548 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$27056 \$153 \$481 \$78 \$273 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27057 \$153 \$606 \$44 \$604 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27059 \$16 \$674 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27061 \$16 \$273 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27062 \$16 \$241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27063 \$153 \$301 \$112 \$115 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27064 \$153 \$481 \$389 \$115 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27065 \$153 \$547 \$559 \$604 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27066 \$153 \$482 \$388 \$115 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27067 \$16 \$354 \$16 \$153 \$115 VNB sky130_fd_sc_hd__inv_1
X$27068 \$153 \$334 \$266 \$485 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27071 \$153 \$363 \$189 \$424 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27072 \$153 \$189 \$591 \$439 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$27073 \$153 \$483 \$389 \$485 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27075 \$153 \$484 \$388 \$485 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27076 \$16 \$151 \$16 \$153 \$485 VNB sky130_fd_sc_hd__inv_1
X$27079 \$16 \$241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27080 \$153 \$364 \$267 \$241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27081 \$153 \$486 \$353 \$177 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27082 \$153 \$576 \$559 \$607 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27083 \$16 \$608 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27085 \$153 \$42 \$559 \$485 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27086 \$16 \$424 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27087 \$153 \$577 \$593 \$424 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27088 \$153 \$577 \$353 \$771 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27090 \$16 \$273 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27092 \$153 \$305 \$81 \$424 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27093 \$16 \$424 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27094 \$16 \$79 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27095 \$153 \$440 \$593 \$79 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27096 \$153 \$488 \$21 \$771 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27097 \$153 \$609 \$44 \$771 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27098 \$16 \$306 \$16 \$153 \$117 VNB sky130_fd_sc_hd__inv_1
X$27102 \$153 \$578 \$425 \$273 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27103 \$153 \$578 \$389 \$348 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27104 \$16 \$441 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27106 \$16 \$79 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27107 \$153 \$366 \$425 \$79 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27110 \$153 \$610 \$559 \$611 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27111 \$16 \$145 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27112 \$153 \$367 \$425 \$145 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27114 \$16 \$508 \$16 \$153 \$348 VNB sky130_fd_sc_hd__inv_1
X$27115 \$153 \$579 \$21 \$348 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27116 \$16 \$723 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27117 \$16 \$508 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27119 \$153 \$83 \$387 \$490 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$27121 \$153 \$391 \$558 \$632 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$27122 \$16 \$387 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27125 \$16 \$509 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27126 \$16 \$446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27127 \$16 \$426 \$16 \$153 \$121 VNB sky130_fd_sc_hd__inv_1
X$27129 \$153 \$633 \$391 \$446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27130 \$153 \$390 \$371 \$121 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27132 \$153 \$524 \$703 \$442 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27133 \$16 \$594 \$16 \$153 \$442 VNB sky130_fd_sc_hd__inv_1
X$27134 \$16 \$149 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27135 \$16 \$63 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27136 \$16 \$178 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27138 \$16 \$310 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27139 \$153 \$525 \$391 \$178 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27140 \$16 \$509 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27142 \$153 \$443 \$391 \$509 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27143 \$16 \$149 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27145 \$153 \$84 \$595 \$634 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$27146 \$153 \$525 \$549 \$442 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27147 \$153 \$550 \$84 \$509 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27149 \$153 \$612 \$57 \$442 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27151 \$153 \$560 \$596 \$149 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27152 \$153 \$368 \$398 \$442 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27154 \$16 \$265 \$428 \$551 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$27155 \$153 \$85 \$423 \$551 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$27158 \$153 \$552 \$85 \$509 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27159 \$16 \$149 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27160 \$16 \$438 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27161 \$153 \$552 \$371 \$122 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27162 \$16 \$438 \$369 \$526 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$27163 \$153 \$427 \$631 \$526 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$27164 \$16 \$369 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27167 \$153 \$400 \$393 \$258 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27168 \$16 \$149 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27169 \$16 \$310 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27170 \$153 \$527 \$427 \$310 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27172 \$16 \$309 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27173 \$153 \$491 \$23 \$502 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27174 \$153 \$492 \$398 \$502 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27175 \$153 \$527 \$223 \$502 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27176 \$153 \$494 \$427 \$178 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27177 \$153 \$493 \$371 \$124 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27179 \$153 \$528 \$427 \$509 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27180 \$153 \$494 \$549 \$502 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27181 \$153 \$528 \$371 \$502 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27182 \$153 \$86 \$591 \$495 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$27183 \$16 \$829 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27184 \$16 \$306 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27186 \$16 \$608 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27187 \$16 \$428 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27188 \$16 \$428 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27189 \$16 \$306 \$428 \$580 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$27190 \$153 \$87 \$116 \$497 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$27191 \$153 \$50 \$608 \$580 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$27192 \$153 \$444 \$87 \$309 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27193 \$16 \$309 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27195 \$16 \$509 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27197 \$153 \$613 \$393 \$445 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27198 \$153 \$373 \$87 \$446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27199 \$16 \$446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27200 \$153 \$510 \$676 \$149 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27201 \$16 \$80 \$16 \$153 \$179 VNB sky130_fd_sc_hd__inv_1
X$27203 \$16 \$509 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27204 \$153 \$614 \$57 \$445 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27207 \$153 \$374 \$50 \$509 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27208 \$16 \$1600 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27209 \$16 \$615 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27210 \$153 \$277 \$1600 \$635 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$27211 \$153 \$510 \$398 \$445 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27213 \$16 \$63 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27214 \$16 \$63 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27216 \$153 \$498 \$277 \$509 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27217 \$153 \$636 \$597 \$63 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27219 \$16 \$306 \$16 \$153 \$126 VNB sky130_fd_sc_hd__inv_1
X$27220 \$153 \$498 \$371 \$181 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27221 \$16 \$615 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27223 \$16 \$178 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27224 \$153 \$581 \$597 \$178 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27227 \$16 \$149 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27228 \$16 \$446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27229 \$153 \$447 \$277 \$446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27230 \$153 \$581 \$549 \$637 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27232 \$16 \$446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27233 \$153 \$499 \$597 \$446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27234 \$16 \$508 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27237 \$153 \$499 \$393 \$637 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27238 \$153 \$638 \$23 \$637 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27239 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$27240 \$153 \$616 \$398 \$637 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27243 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$27244 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$27245 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$27246 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$27247 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$27248 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$27249 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$27250 \$153 \$2582 \$2510 \$1687 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27251 \$153 \$2470 \$2510 \$2006 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27252 \$16 \$1687 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27254 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$27255 \$153 \$2470 \$1943 \$2343 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27259 \$153 \$2351 \$2510 \$1795 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27260 \$153 \$2532 \$2510 \$1942 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27261 \$153 \$2583 \$2510 \$2024 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27262 \$16 \$1942 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27263 \$16 \$1795 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27264 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$27266 \$153 \$2471 \$2510 \$2180 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27267 \$16 \$2024 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27268 \$16 \$1037 \$16 \$153 \$2343 VNB sky130_fd_sc_hd__inv_1
X$27270 \$153 \$2440 \$2377 \$1687 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27271 \$153 \$2471 \$2252 \$2343 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27272 \$16 \$2180 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27273 \$16 \$1658 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27275 \$16 \$2006 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27276 \$153 \$2583 \$2210 \$2343 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27277 \$153 \$2472 \$2377 \$2006 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27278 \$153 \$2574 \$2210 \$2110 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27279 \$153 \$2472 \$1943 \$2179 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27280 \$16 \$1687 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27281 \$16 \$1291 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27282 \$153 \$2584 \$2511 \$2180 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27284 \$153 \$2497 \$2064 \$2179 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27286 \$16 \$2180 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27287 \$153 \$2249 \$2511 \$1795 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27289 \$153 \$2473 \$2511 \$1687 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27290 \$16 \$2006 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27292 \$16 \$1013 \$16 \$153 \$2275 VNB sky130_fd_sc_hd__inv_1
X$27293 \$153 \$2441 \$2064 \$1861 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27294 \$153 \$2511 \$972 \$2512 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$27295 \$16 \$1013 \$1522 \$2512 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$27296 \$153 \$2575 \$2380 \$2006 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27297 \$153 \$2137 \$2009 \$1861 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27300 \$153 \$2533 \$2380 \$1687 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27301 \$153 \$2473 \$1792 \$2275 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27302 \$153 \$2620 \$2064 \$2275 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27304 \$16 \$2006 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27305 \$16 \$1067 \$1522 \$2534 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$27307 \$16 \$1348 \$2932 \$2585 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$27308 \$153 \$2474 \$2354 \$2006 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27309 \$16 \$1980 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27311 \$153 \$2250 \$2354 \$1942 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27312 \$153 \$2474 \$1943 \$2181 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27313 \$16 \$1942 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27314 \$16 \$2932 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27315 \$153 \$2551 \$2354 \$2024 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27316 \$16 \$1522 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27318 \$16 \$1522 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27319 \$16 \$1980 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27321 \$153 \$2417 \$2354 \$2180 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27322 \$153 \$2587 \$2009 \$2586 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27323 \$16 \$2180 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27324 \$153 \$2551 \$2210 \$2181 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27326 \$153 \$2475 \$2290 \$1980 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27327 \$16 \$2024 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27329 \$16 \$2442 \$16 \$153 \$1522 VNB sky130_fd_sc_hd__clkbuf_2
X$27330 \$16 \$1795 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27331 \$153 \$2588 \$2210 \$2344 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27333 \$153 \$2443 \$2252 \$2344 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27335 \$16 \$2180 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27336 \$153 \$2475 \$2009 \$2344 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27338 \$153 \$2552 \$2290 \$1795 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27339 \$16 \$2006 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27341 \$153 \$2476 \$2290 \$2006 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27342 \$153 \$2552 \$1815 \$2344 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27343 \$153 \$2476 \$1943 \$2344 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27344 \$16 \$1942 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27346 \$153 \$2535 \$1815 \$2386 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27348 \$153 \$2535 \$2478 \$1795 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27351 \$153 \$2589 \$2478 \$1687 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27352 \$153 \$2385 \$2064 \$2219 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27353 \$16 \$1687 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27354 \$16 \$1795 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27355 \$16 \$2647 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27357 \$16 \$2479 \$16 \$153 \$1048 VNB sky130_fd_sc_hd__clkbuf_2
X$27358 \$16 \$2006 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27359 \$153 \$2553 \$2478 \$2006 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27361 \$153 \$2477 \$2478 \$2180 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27362 \$153 \$2553 \$1943 \$2386 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27363 \$16 \$2113 \$16 \$153 \$2436 VNB sky130_fd_sc_hd__clkbuf_2
X$27364 \$153 \$2536 \$2478 \$1658 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27365 \$16 \$1048 \$2647 \$2590 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$27368 \$16 \$2100 \$16 \$153 \$2434 VNB sky130_fd_sc_hd__clkbuf_2
X$27369 \$153 \$2536 \$1547 \$2386 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27370 \$153 \$2537 \$2478 \$1980 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27371 \$153 \$2591 \$1815 \$2634 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27372 \$16 \$2576 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27373 \$16 \$2576 \$16 \$153 \$2113 VNB sky130_fd_sc_hd__clkbuf_2
X$27374 \$153 \$2479 \$2436 \$2435 \$2434 \$2420 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$27376 \$153 \$2513 \$2434 \$2435 \$2436 \$2420 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$27377 \$16 \$2936 \$16 \$153 \$2195 VNB sky130_fd_sc_hd__clkbuf_2
X$27378 \$16 \$2936 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27379 \$16 \$1980 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27382 \$153 \$2436 \$2434 \$2355 \$2420 \$2435 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$27383 \$153 \$2436 \$2420 \$2356 \$2434 \$2435 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$27384 \$153 \$2434 \$2420 \$2480 \$2436 \$2435 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$27385 \$16 \$1037 \$2539 \$2592 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$27388 \$16 \$2294 \$16 \$153 \$2538 VNB sky130_fd_sc_hd__clkbuf_2
X$27389 \$16 \$2539 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27391 \$153 \$2421 \$2389 \$2199 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27392 \$153 \$2481 \$2389 \$1965 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27393 \$153 \$2577 \$2184 \$2594 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27394 \$16 \$2513 \$16 \$153 \$1264 VNB sky130_fd_sc_hd__clkbuf_2
X$27395 \$16 \$1965 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27397 \$153 \$2447 \$2389 \$2089 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27398 \$16 \$2480 \$16 \$153 \$588 VNB sky130_fd_sc_hd__clkbuf_2
X$27399 \$16 \$2199 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27400 \$153 \$2446 \$1924 \$2390 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27401 \$153 \$2593 \$1924 \$2594 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27402 \$16 \$2514 \$16 \$153 \$1508 VNB sky130_fd_sc_hd__clkbuf_2
X$27404 \$153 \$2357 \$2389 \$2043 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27405 \$16 \$2089 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27408 \$153 \$2391 \$2389 \$1805 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27409 \$16 \$2043 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27410 \$153 \$2498 \$1471 \$2594 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27411 \$16 \$1805 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27413 \$16 \$1553 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27414 \$16 \$1805 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27415 \$153 \$2595 \$2244 \$2043 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27416 \$16 \$1348 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27417 \$16 \$972 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27418 \$16 \$2539 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27420 \$153 \$2448 \$2244 \$2089 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27421 \$16 \$2043 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27423 \$16 \$2089 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27424 \$153 \$2555 \$972 \$2554 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$27425 \$16 \$2089 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27426 \$153 \$2540 \$2244 \$2199 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27429 \$153 \$2540 \$2184 \$2299 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27430 \$153 \$2406 \$1924 \$2299 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27431 \$153 \$2556 \$2555 \$2089 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27432 \$153 \$2393 \$1895 \$2299 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27433 \$16 \$2199 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27434 \$16 \$2199 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27435 \$16 \$1013 \$16 \$153 \$2557 VNB sky130_fd_sc_hd__inv_1
X$27437 \$153 \$2449 \$2184 \$1922 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27438 \$16 \$2089 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27439 \$153 \$2558 \$2555 \$2042 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27440 \$16 \$1013 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27441 \$16 \$1291 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27442 \$16 \$1845 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27443 \$153 \$2515 \$2184 \$2327 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27444 \$153 \$2625 \$1471 \$2557 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27445 \$153 \$2361 \$2359 \$2042 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27447 \$153 \$2515 \$2359 \$2199 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27448 \$16 \$2042 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27449 \$153 \$2525 \$1211 \$2451 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$27450 \$16 \$2199 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27451 \$16 \$1047 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27452 \$16 \$1211 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27454 \$153 \$2559 \$2525 \$1845 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27457 \$16 \$1845 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27458 \$16 \$1067 \$16 \$153 \$2499 VNB sky130_fd_sc_hd__inv_1
X$27459 \$153 \$2482 \$2525 \$1805 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27460 \$153 \$2452 \$2525 \$2199 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27462 \$153 \$2482 \$1703 \$2499 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27465 \$153 \$2597 \$842 \$2596 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$27466 \$16 \$2362 \$16 \$153 \$2347 VNB sky130_fd_sc_hd__clkbuf_2
X$27467 \$16 \$1805 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27468 \$16 \$842 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27469 \$153 \$2541 \$2277 \$1805 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27470 \$153 \$2526 \$2277 \$2089 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27472 \$16 \$1805 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27473 \$153 \$2541 \$1703 \$2152 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27474 \$153 \$2526 \$2026 \$2152 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27475 \$16 \$1048 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27476 \$16 \$2089 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27477 \$16 \$1048 \$2347 \$2542 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$27479 \$153 \$2560 \$1173 \$2542 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$27480 \$153 \$2453 \$2200 \$2199 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27482 \$16 \$1173 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27483 \$153 \$2598 \$1471 \$2186 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27484 \$16 \$2199 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27485 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$27486 \$153 \$2543 \$2200 \$2043 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27487 \$153 \$2454 \$2200 \$1805 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27488 \$153 \$2543 \$1954 \$2186 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27490 \$16 \$2043 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27491 \$16 \$1805 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27492 \$16 \$584 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27495 \$153 \$2483 \$2365 \$2042 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27496 \$153 \$2527 \$2365 \$2199 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27497 \$153 \$2483 \$1924 \$2120 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27498 \$16 \$2042 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27501 \$153 \$2599 \$2578 \$1923 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27502 \$153 \$2527 \$2184 \$2120 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27503 \$16 \$716 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27505 \$16 \$2043 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27506 \$153 \$2516 \$1703 \$2500 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27507 \$153 \$2528 \$2365 \$2043 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27510 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$27511 \$16 \$2089 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27512 \$153 \$2600 \$2578 \$2089 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27513 \$153 \$2528 \$1954 \$2120 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27514 \$153 \$2455 \$1471 \$2120 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27515 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$27517 \$153 \$2303 \$2517 \$1879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27519 \$153 \$2601 \$2517 \$2098 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27520 \$153 \$2456 \$1558 \$2278 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27521 \$16 \$2098 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27523 \$16 \$902 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27524 \$16 \$1459 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27525 \$16 \$1879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27526 \$16 \$3272 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27527 \$153 \$2602 \$2517 \$1878 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27528 \$16 \$1756 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27530 \$153 \$2484 \$2279 \$1756 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27531 \$153 \$2517 \$1459 \$2603 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$27532 \$153 \$2484 \$1712 \$2278 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27534 \$16 \$902 \$16 \$153 \$2161 VNB sky130_fd_sc_hd__inv_1
X$27535 \$16 \$2104 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27537 \$153 \$2501 \$2485 \$2105 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27538 \$153 \$2561 \$2485 \$2104 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27540 \$153 \$2501 \$2438 \$2502 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27541 \$153 \$2561 \$2092 \$2502 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27543 \$16 \$2105 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27544 \$16 \$1756 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27547 \$153 \$2544 \$2485 \$1756 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27548 \$153 \$2562 \$2485 \$1879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27550 \$153 \$2544 \$1712 \$2502 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27551 \$16 \$438 \$16 \$153 \$2502 VNB sky130_fd_sc_hd__inv_1
X$27552 \$153 \$2485 \$631 \$2457 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$27553 \$16 \$595 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27555 \$16 \$1543 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27557 \$16 \$2105 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27558 \$153 \$1827 \$353 \$1811 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27559 \$16 \$631 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27561 \$16 \$2098 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27562 \$153 \$2486 \$2202 \$2098 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27563 \$153 \$2503 \$2202 \$2105 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27566 \$153 \$2486 \$1993 \$2280 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27567 \$16 \$1245 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27568 \$16 \$1933 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27569 \$16 \$2104 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27570 \$153 \$2604 \$2202 \$2104 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27571 \$153 \$2503 \$2438 \$2280 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27573 \$16 \$1456 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27574 \$153 \$2458 \$1868 \$2280 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27575 \$16 \$2232 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27576 \$16 \$1585 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27578 \$16 \$2098 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27579 \$153 \$2487 \$2309 \$2105 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27580 \$16 \$2104 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27581 \$153 \$2563 \$2309 \$2104 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27583 \$153 \$2487 \$2438 \$2334 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27584 \$153 \$2563 \$2092 \$2334 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27587 \$153 \$2460 \$2309 \$2016 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27588 \$153 \$2459 \$1558 \$2334 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27589 \$16 \$1969 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27590 \$153 \$2564 \$2579 \$1969 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27591 \$16 \$2016 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27593 \$16 \$2016 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27594 \$153 \$2399 \$2310 \$2016 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27596 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$27598 \$153 \$2605 \$1993 \$2606 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27599 \$16 \$2105 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27600 \$153 \$2488 \$2310 \$2105 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27601 \$153 \$2564 \$1613 \$2606 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27603 \$16 \$2580 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27605 \$153 \$2488 \$2438 \$2187 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27606 \$153 \$2607 \$1715 \$2606 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27607 \$153 \$2425 \$2092 \$2187 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27608 \$16 \$1879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27609 \$16 \$1184 \$2580 \$2608 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$27610 \$153 \$2565 \$2092 \$2606 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27611 \$153 \$2461 \$1558 \$2187 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27613 \$16 \$1756 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27614 \$16 \$2104 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27616 \$153 \$2489 \$2368 \$2104 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27617 \$153 \$2609 \$2368 \$1756 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27618 \$153 \$2489 \$2092 \$2188 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27620 \$16 \$1969 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27621 \$153 \$2566 \$2732 \$1969 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27622 \$16 \$1811 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27624 \$16 \$1879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27625 \$153 \$2490 \$2368 \$1879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27627 \$16 \$1445 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27628 \$153 \$2843 \$1558 \$2504 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27629 \$153 \$2490 \$1558 \$2188 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27630 \$153 \$2566 \$1613 \$2504 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27631 \$16 \$2105 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27633 \$16 \$508 \$2580 \$2545 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$27634 \$153 \$2518 \$2732 \$2105 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27635 \$153 \$2518 \$2438 \$2504 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27636 \$16 \$276 \$16 \$153 \$2504 VNB sky130_fd_sc_hd__inv_1
X$27637 \$16 \$723 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27638 \$16 \$276 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27639 \$16 \$2314 \$16 \$153 \$2733 VNB sky130_fd_sc_hd__clkbuf_2
X$27640 \$16 \$508 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27641 \$16 \$895 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27642 \$16 \$2189 \$16 \$153 \$2337 VNB sky130_fd_sc_hd__clkbuf_2
X$27643 \$16 \$2519 \$16 \$153 \$1518 VNB sky130_fd_sc_hd__clkbuf_2
X$27644 \$16 \$2204 \$16 \$153 \$2371 VNB sky130_fd_sc_hd__clkbuf_2
X$27647 \$153 \$2520 \$2371 \$2464 \$2372 \$2337 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$27648 \$16 \$2520 \$16 \$153 \$2462 VNB sky130_fd_sc_hd__clkbuf_2
X$27649 \$16 \$2521 \$16 \$153 \$1120 VNB sky130_fd_sc_hd__clkbuf_2
X$27650 \$16 \$2505 \$16 \$153 \$1184 VNB sky130_fd_sc_hd__clkbuf_2
X$27651 \$153 \$2521 \$2372 \$2464 \$2371 \$2337 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$27652 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$27653 \$153 \$2372 \$2371 \$2465 \$2337 \$2464 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$27655 \$16 \$902 \$1972 \$2610 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$27656 \$16 \$2464 \$2337 \$2372 \$2371 \$16 \$153 \$2734 VNB
+ sky130_fd_sc_hd__and4_2
X$27658 \$153 \$2612 \$1459 \$2610 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$27660 \$153 \$2547 \$2316 \$2085 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27661 \$16 \$2611 \$16 \$153 \$508 VNB sky130_fd_sc_hd__clkbuf_2
X$27662 \$16 \$1459 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27663 \$153 \$2547 \$2271 \$2402 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27664 \$16 \$2085 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27665 \$16 \$594 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27667 \$16 \$2031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27668 \$16 \$902 \$16 \$153 \$2613 VNB sky130_fd_sc_hd__inv_1
X$27669 \$16 \$902 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27670 \$153 \$2522 \$2056 \$2402 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27671 \$153 \$2522 \$2316 \$1973 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27672 \$153 \$2548 \$2316 \$1860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27673 \$16 \$1973 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27674 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$27676 \$153 \$2548 \$2000 \$2402 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27677 \$16 \$1860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27678 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$27679 \$16 \$2232 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27680 \$153 \$2549 \$1935 \$2192 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27682 \$153 \$2567 \$1935 \$1860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27683 \$16 \$2192 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27684 \$16 \$2031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27685 \$153 \$2549 \$2269 \$2506 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27687 \$16 \$1860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27688 \$16 \$2093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27689 \$153 \$2492 \$1935 \$2031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27690 \$153 \$2567 \$2000 \$2506 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27692 \$16 \$631 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27693 \$153 \$2614 \$2056 \$2506 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27694 \$153 \$2581 \$631 \$2467 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$27696 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$27697 \$16 \$1960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27699 \$153 \$2568 \$2581 \$1960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27700 \$153 \$2237 \$1936 \$1870 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27701 \$153 \$2529 \$2271 \$2506 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27702 \$153 \$2568 \$2086 \$2491 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27703 \$16 \$438 \$16 \$153 \$2491 VNB sky130_fd_sc_hd__inv_1
X$27705 \$153 \$2507 \$2000 \$2491 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27706 \$16 \$438 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27708 \$16 \$2093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27709 \$153 \$2569 \$2581 \$2093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27710 \$153 \$2492 \$1936 \$2506 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27712 \$153 \$2781 \$2271 \$2491 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27714 \$16 \$1719 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27716 \$153 \$2569 \$2265 \$2491 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27717 \$153 \$2834 \$2056 \$2780 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27718 \$16 \$1184 \$2531 \$2550 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$27720 \$153 \$2530 \$2570 \$2031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27721 \$16 \$2031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27722 \$16 \$1184 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27723 \$16 \$1514 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27724 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$27725 \$16 \$1184 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27726 \$16 \$1860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27727 \$16 \$1184 \$16 \$153 \$2508 VNB sky130_fd_sc_hd__inv_1
X$27729 \$153 \$2530 \$1936 \$2508 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27730 \$153 \$2571 \$2570 \$1860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27731 \$153 \$2468 \$2265 \$2239 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27732 \$153 \$2571 \$2000 \$2508 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27734 \$16 \$508 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27735 \$16 \$1973 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27736 \$153 \$2493 \$2403 \$1973 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27737 \$16 \$2192 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27739 \$153 \$2615 \$2403 \$2192 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27741 \$153 \$2469 \$2000 \$2282 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27743 \$16 \$508 \$2531 \$2616 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$27744 \$16 \$2191 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27745 \$16 \$724 \$2531 \$2494 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$27746 \$153 \$2523 \$2403 \$2191 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27748 \$16 \$2031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27749 \$153 \$2523 \$2267 \$2282 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27750 \$16 \$276 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27751 \$153 \$2524 \$895 \$2494 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$27752 \$153 \$2572 \$723 \$2616 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$27753 \$153 \$2495 \$2524 \$2085 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27754 \$16 \$2191 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27756 \$153 \$2573 \$2267 \$2032 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27757 \$153 \$2573 \$2524 \$2191 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27758 \$16 \$724 \$16 \$153 \$2032 VNB sky130_fd_sc_hd__inv_1
X$27759 \$16 \$276 \$16 \$153 \$2284 VNB sky130_fd_sc_hd__inv_1
X$27760 \$153 \$2509 \$2000 \$2178 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27762 \$16 \$1860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27765 \$153 \$2496 \$2524 \$1860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27766 \$16 \$2031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27767 \$153 \$2617 \$2269 \$2178 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27768 \$153 \$2063 \$2524 \$2031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27769 \$153 \$2131 \$2524 \$1973 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27772 \$16 \$2192 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27773 \$153 \$2132 \$2524 \$2192 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27774 \$153 \$2207 \$2524 \$1960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27775 \$153 \$2618 \$2269 \$2642 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27776 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$27778 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$27779 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$27780 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$27781 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$27782 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$27783 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$27784 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$27785 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$27788 \$153 \$1494 \$1256 \$263 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27789 \$153 \$1388 \$1256 \$17 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27790 \$153 \$1388 \$102 \$1187 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27792 \$16 \$504 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27793 \$16 \$263 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27795 \$16 \$17 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27798 \$153 \$1495 \$1465 \$395 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27799 \$153 \$1427 \$1256 \$395 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27800 \$16 \$395 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27801 \$16 \$395 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27802 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$27804 \$16 \$1496 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27806 \$16 \$1168 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27808 \$153 \$1497 \$1465 \$419 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27809 \$16 \$783 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27810 \$16 \$1390 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27811 \$153 \$1428 \$1256 \$184 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27812 \$153 \$1495 \$394 \$1535 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27813 \$153 \$1428 \$59 \$1187 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27814 \$16 \$1496 \$16 \$153 \$1535 VNB sky130_fd_sc_hd__inv_1
X$27816 \$16 \$419 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27817 \$16 \$184 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27818 \$16 \$1496 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27819 \$153 \$1450 \$1257 \$419 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27820 \$153 \$1429 \$1257 \$504 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27821 \$153 \$1450 \$349 \$1106 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27822 \$16 \$419 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27823 \$16 \$504 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27825 \$16 \$1430 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27826 \$16 \$1480 \$16 \$153 \$1106 VNB sky130_fd_sc_hd__inv_1
X$27829 \$16 \$1480 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27830 \$16 \$1168 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27831 \$16 \$1404 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27832 \$153 \$1451 \$1326 \$419 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27833 \$153 \$1431 \$1326 \$17 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27834 \$16 \$1404 \$1168 \$1498 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$27835 \$16 \$249 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27836 \$16 \$504 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27837 \$16 \$419 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27838 \$153 \$1432 \$1326 \$395 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27841 \$153 \$1417 \$1326 \$263 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27842 \$153 \$1432 \$394 \$1327 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27843 \$16 \$263 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27844 \$16 \$504 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27845 \$153 \$1418 \$1249 \$504 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27846 \$16 \$395 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27847 \$16 \$58 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27848 \$16 \$1404 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27850 \$153 \$1417 \$234 \$1327 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27852 \$153 \$1499 \$1249 \$249 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27853 \$153 \$1346 \$349 \$1250 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27854 \$153 \$1418 \$561 \$1250 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27855 \$16 \$1328 \$16 \$153 \$1250 VNB sky130_fd_sc_hd__inv_1
X$27856 \$153 \$1347 \$234 \$1250 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27858 \$16 \$249 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27859 \$16 \$395 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27860 \$16 \$263 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27861 \$16 \$419 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27862 \$153 \$1405 \$1258 \$249 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27863 \$153 \$1329 \$1258 \$419 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27864 \$16 \$249 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27865 \$153 \$1500 \$1258 \$263 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27866 \$16 \$1433 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27868 \$153 \$1405 \$377 \$1191 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27869 \$16 \$1433 \$16 \$153 \$1192 VNB sky130_fd_sc_hd__clkbuf_2
X$27870 \$153 \$1501 \$1330 \$249 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27871 \$153 \$1434 \$1330 \$504 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27874 \$153 \$1210 \$234 \$1193 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27875 \$153 \$1284 \$349 \$1193 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27877 \$16 \$504 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27878 \$153 \$1453 \$1330 \$419 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27880 \$153 \$1330 \$1139 \$1350 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$27881 \$153 \$1453 \$349 \$1454 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27883 \$16 \$1264 \$715 \$1351 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$27884 \$153 \$1435 \$1352 \$17 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27885 \$16 \$419 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27887 \$153 \$1481 \$349 \$1251 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27888 \$153 \$1435 \$102 \$1251 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27889 \$16 \$395 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27890 \$16 \$1264 \$16 \$153 \$1251 VNB sky130_fd_sc_hd__inv_1
X$27891 \$153 \$1389 \$1352 \$395 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27893 \$153 \$1466 \$377 \$1251 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27895 \$153 \$1467 \$59 \$1251 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27896 \$153 \$1353 \$561 \$1251 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27897 \$153 \$1349 \$234 \$1454 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27898 \$16 \$504 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27899 \$16 \$1331 \$430 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$27901 \$153 \$1068 \$349 \$1070 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27902 \$153 \$1406 \$504 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$27903 \$153 \$1155 \$394 \$1070 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27904 \$153 \$1127 \$234 \$1070 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27905 \$16 \$1406 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27906 \$153 \$1407 \$395 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$27909 \$16 \$1482 \$16 \$153 \$1502 VNB sky130_fd_sc_hd__clkbuf_2
X$27910 \$16 \$1502 \$16 \$153 \$1182 VNB sky130_fd_sc_hd__clkbuf_2
X$27911 \$16 \$1331 \$1263 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$27912 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27913 \$16 \$1331 \$1211 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$27914 \$153 \$153 \$30 \$1408 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27915 \$16 \$1436 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27916 \$153 \$153 \$377 \$1408 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27917 \$153 \$153 \$349 \$1408 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27919 \$153 \$153 \$59 \$1408 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27920 \$153 \$153 \$394 \$1408 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27921 \$153 \$153 \$102 \$1408 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27922 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27923 \$153 \$1261 \$1503 \$1468 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$27924 \$16 \$1390 \$979 \$1355 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$27925 \$16 \$394 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27927 \$153 \$1437 \$1261 \$187 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27929 \$16 \$1496 \$979 \$1468 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$27930 \$16 \$979 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27931 \$16 \$979 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27932 \$16 \$979 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27933 \$16 \$1390 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27934 \$16 \$1496 \$16 \$153 \$1409 VNB sky130_fd_sc_hd__inv_1
X$27935 \$153 \$1437 \$54 \$1409 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27936 \$153 \$1308 \$346 \$1409 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27937 \$153 \$1505 \$1504 \$358 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27938 \$16 \$1390 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27940 \$16 \$1496 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27941 \$16 \$1332 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27942 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$27943 \$153 \$1356 \$215 \$1409 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27944 \$16 \$358 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27945 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$27946 \$153 \$1469 \$253 \$1409 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27947 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$27949 \$153 \$1438 \$1261 \$212 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27950 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$27952 \$153 \$1506 \$1504 \$18 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27953 \$153 \$1357 \$104 \$1409 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27954 \$153 \$1438 \$347 \$1409 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27955 \$16 \$212 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27956 \$16 \$981 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27957 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$27958 \$16 \$18 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27961 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$27962 \$153 \$1289 \$35 \$1333 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27963 \$153 \$1391 \$1262 \$358 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27964 \$153 \$1470 \$346 \$1333 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27965 \$153 \$1507 \$1471 \$1483 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27966 \$153 \$1392 \$1262 \$60 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27969 \$153 \$1484 \$347 \$1333 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27970 \$153 \$1392 \$104 \$1333 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27971 \$16 \$60 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27972 \$16 \$753 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27974 \$16 \$710 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27975 \$153 \$1419 \$1334 \$60 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27976 \$16 \$1292 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27978 \$16 \$1291 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27979 \$153 \$1419 \$104 \$1393 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27980 \$153 \$1358 \$215 \$1393 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27981 \$153 \$1359 \$1334 \$358 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27982 \$16 \$60 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27983 \$16 \$1328 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27984 \$16 \$18 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27985 \$153 \$1158 \$347 \$1040 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27986 \$153 \$1394 \$1334 \$18 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27988 \$153 \$1528 \$54 \$1393 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27989 \$16 \$187 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27990 \$153 \$1420 \$1421 \$358 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27991 \$16 \$293 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27992 \$16 \$358 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27994 \$16 \$1485 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$27995 \$153 \$1420 \$253 \$1335 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$27996 \$16 \$1485 \$16 \$153 \$908 VNB sky130_fd_sc_hd__clkbuf_2
X$27997 \$153 \$1360 \$1421 \$73 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$27999 \$153 \$1439 \$1421 \$60 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28000 \$16 \$908 \$16 \$153 \$946 VNB sky130_fd_sc_hd__clkbuf_2
X$28002 \$16 \$60 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28003 \$16 \$691 \$946 \$1440 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$28005 \$153 \$1472 \$842 \$1440 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$28006 \$153 \$1041 \$1171 \$1395 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$28007 \$16 \$18 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28008 \$153 \$1159 \$35 \$1040 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28009 \$16 \$691 \$16 \$153 \$1410 VNB sky130_fd_sc_hd__inv_1
X$28010 \$153 \$1441 \$1472 \$18 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28011 \$16 \$358 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28014 \$153 \$1361 \$253 \$1199 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28015 \$16 \$18 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28016 \$153 \$1422 \$1472 \$358 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28017 \$153 \$1362 \$346 \$1199 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28018 \$16 \$351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28019 \$153 \$1422 \$253 \$1410 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28020 \$16 \$358 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28023 \$16 \$1171 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28024 \$153 \$911 \$1336 \$18 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28025 \$16 \$1264 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28026 \$16 \$1173 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28027 \$16 \$1048 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28028 \$153 \$1486 \$54 \$1410 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28029 \$16 \$1508 \$16 \$153 \$1411 VNB sky130_fd_sc_hd__inv_1
X$28030 \$153 \$1423 \$1336 \$187 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28033 \$153 \$1442 \$1336 \$212 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28034 \$153 \$1442 \$347 \$1411 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28035 \$153 \$1423 \$54 \$1411 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28036 \$16 \$187 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28037 \$153 \$153 \$253 \$1487 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28038 \$16 \$212 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28039 \$153 \$1200 \$1336 \$73 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28041 \$153 \$153 \$104 \$1487 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28042 \$16 \$16 \$153 VNB sky130_fd_sc_hd__conb_1
X$28044 \$153 \$1488 \$73 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$28045 \$153 \$1366 \$104 \$1411 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28046 \$16 \$73 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28047 \$16 \$1407 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28050 \$153 \$1367 \$358 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$28051 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28055 \$16 \$1436 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28056 \$153 \$1474 \$44 \$1811 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28057 \$153 \$1436 \$145 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$28058 \$153 \$1132 \$388 \$947 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28059 \$16 \$1543 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28060 \$16 \$1446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28061 \$16 \$399 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28064 \$153 \$153 \$21 \$1337 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28065 \$16 \$559 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28066 \$16 \$1378 \$16 \$153 \$1337 VNB sky130_fd_sc_hd__clkbuf_2
X$28067 \$153 \$153 \$388 \$1337 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28068 \$153 \$153 \$266 \$1337 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28069 \$153 \$153 \$112 \$1337 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28070 \$153 \$153 \$44 \$1337 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28071 \$16 \$145 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28073 \$153 \$1509 \$1183 \$273 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28074 \$153 \$1443 \$1183 \$145 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28075 \$153 \$408 \$21 \$604 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28078 \$16 \$1929 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28079 \$16 \$273 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28080 \$16 \$145 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28081 \$16 \$82 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28082 \$153 \$1444 \$1268 \$145 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28083 \$153 \$1511 \$1268 \$273 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28084 \$16 \$1566 \$1446 \$1512 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$28085 \$153 \$1225 \$112 \$657 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28088 \$153 \$1510 \$21 \$1252 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28089 \$153 \$1318 \$559 \$1252 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28091 \$16 \$82 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28092 \$153 \$1445 \$1338 \$79 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28093 \$153 \$1474 \$1338 \$82 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28095 \$153 \$1238 \$559 \$1396 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28096 \$153 \$1455 \$1338 \$145 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28097 \$153 \$1298 \$112 \$1396 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28098 \$16 \$145 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28099 \$16 \$1201 \$16 \$153 \$1446 VNB sky130_fd_sc_hd__clkbuf_2
X$28101 \$153 \$1447 \$44 \$1541 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28102 \$153 \$1447 \$1253 \$82 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28104 \$153 \$1513 \$1253 \$145 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28105 \$153 \$722 \$21 \$913 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28106 \$16 \$145 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28107 \$153 \$937 \$266 \$913 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28108 \$16 \$1446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28109 \$16 \$1566 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28111 \$153 \$742 \$112 \$913 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28114 \$153 \$1598 \$1270 \$82 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28116 \$16 \$441 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28117 \$16 \$1514 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28118 \$16 \$1456 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28119 \$153 \$1397 \$21 \$1412 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28120 \$16 \$1456 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28121 \$16 \$2462 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28124 \$16 \$273 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28125 \$153 \$1371 \$559 \$1412 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28126 \$16 \$82 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28127 \$153 \$1457 \$1254 \$273 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28129 \$16 \$1456 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28130 \$153 \$1457 \$389 \$1412 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28134 \$153 \$1372 \$112 \$1240 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28135 \$16 \$1475 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28136 \$16 \$1184 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28137 \$16 \$145 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28138 \$153 \$1373 \$1320 \$145 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28141 \$153 \$1476 \$389 \$1240 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28142 \$16 \$82 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28143 \$153 \$1476 \$1320 \$273 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28144 \$16 \$273 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28145 \$16 \$424 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28146 \$16 \$441 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28147 \$16 \$82 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28149 \$153 \$1515 \$1424 \$82 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28151 \$16 \$424 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28152 \$153 \$1376 \$559 \$1205 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28153 \$16 \$79 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28154 \$153 \$1398 \$1424 \$79 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28157 \$16 \$1184 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28158 \$16 \$724 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28159 \$16 \$145 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28160 \$153 \$1458 \$1424 \$145 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28162 \$153 \$1413 \$21 \$1229 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28163 \$153 \$1377 \$21 \$1205 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28164 \$153 \$1458 \$266 \$1229 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28166 \$16 \$1367 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28167 \$16 \$1488 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28170 \$153 \$1488 \$310 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$28171 \$153 \$1367 \$309 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$28172 \$16 \$1044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28173 \$16 \$1378 \$16 \$153 \$1243 VNB sky130_fd_sc_hd__clkbuf_2
X$28174 \$16 \$1459 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28177 \$16 \$1489 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28178 \$153 \$153 \$223 \$1243 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28179 \$16 \$1516 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28180 \$153 \$153 \$398 \$1243 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28181 \$153 \$153 \$57 \$1243 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28183 \$153 \$1516 \$149 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$28184 \$16 \$1044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28185 \$16 \$1760 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28186 \$16 \$998 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28187 \$16 \$149 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28189 \$153 \$1449 \$1340 \$149 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28190 \$153 \$1460 \$1340 \$446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28191 \$16 \$595 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28192 \$16 \$399 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28193 \$16 \$310 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28194 \$153 \$1399 \$1340 \$310 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28195 \$16 \$595 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28196 \$16 \$509 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28198 \$153 \$1460 \$393 \$1341 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28199 \$16 \$309 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28200 \$153 \$1399 \$223 \$1341 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28202 \$16 \$310 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28203 \$153 \$1461 \$1565 \$310 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28204 \$153 \$1449 \$398 \$1341 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28206 \$153 \$1277 \$1147 \$178 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28207 \$153 \$1461 \$223 \$1651 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28209 \$16 \$63 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28210 \$153 \$1400 \$1147 \$63 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28211 \$16 \$63 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28213 \$153 \$1490 \$57 \$1651 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28215 \$153 \$748 \$703 \$659 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28216 \$153 \$1400 \$57 \$1059 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28217 \$153 \$1517 \$1622 \$310 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28218 \$153 \$862 \$371 \$659 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28219 \$16 \$1485 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28220 \$16 \$446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28221 \$153 \$1462 \$1622 \$309 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28223 \$153 \$1380 \$393 \$1115 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28224 \$153 \$1401 \$1278 \$63 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28225 \$153 \$1004 \$398 \$659 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28226 \$16 \$63 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28227 \$16 \$1518 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28228 \$153 \$1401 \$57 \$1115 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28232 \$16 \$63 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28233 \$153 \$1519 \$1342 \$63 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28234 \$16 \$149 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28235 \$153 \$1279 \$1342 \$149 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28236 \$153 \$1477 \$398 \$1491 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28237 \$16 \$310 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28239 \$153 \$1478 \$223 \$1255 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28240 \$153 \$1381 \$23 \$1255 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28243 \$16 \$310 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28244 \$16 \$63 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28245 \$153 \$1463 \$1302 \$63 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28248 \$153 \$1382 \$223 \$1343 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28249 \$153 \$1463 \$57 \$1343 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28251 \$16 \$309 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28252 \$153 \$1425 \$1492 \$309 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28253 \$16 \$1514 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28254 \$153 \$1425 \$703 \$1414 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28256 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$28258 \$153 \$1384 \$57 \$776 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28259 \$16 \$1475 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28260 \$16 \$310 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28261 \$153 \$1426 \$1492 \$310 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28262 \$153 \$1385 \$371 \$776 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28264 \$153 \$1426 \$223 \$1414 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28265 \$16 \$1228 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28266 \$16 \$615 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28267 \$16 \$309 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28270 \$16 \$63 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28271 \$16 \$63 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28272 \$153 \$1402 \$1416 \$63 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28273 \$153 \$1464 \$1416 \$309 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28274 \$153 \$1402 \$57 \$1415 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28275 \$153 \$1493 \$398 \$1414 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28277 \$153 \$1464 \$703 \$1415 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28278 \$153 \$1479 \$1416 \$149 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28279 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$28280 \$153 \$1479 \$398 \$1415 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28281 \$16 \$149 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28282 \$16 \$310 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28283 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$28284 \$16 \$310 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28286 \$153 \$1345 \$1416 \$310 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28287 \$153 \$1307 \$393 \$1206 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28288 \$153 \$1403 \$23 \$1415 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28289 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$28292 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$28293 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$28294 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$28295 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$28296 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$28297 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$28298 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$28299 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$28300 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$28301 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$28302 \$153 \$12986 \$13063 \$12230 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28305 \$153 \$13112 \$13063 \$12294 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28307 \$16 \$12294 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28308 \$153 \$13112 \$12208 \$12982 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28309 \$153 \$13044 \$13063 \$12236 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28310 \$16 \$12294 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28311 \$16 \$12230 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28312 \$16 \$11289 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28313 \$16 \$12236 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28315 \$16 \$11289 \$16 \$153 \$12982 VNB sky130_fd_sc_hd__inv_1
X$28316 \$153 \$13129 \$13063 \$12095 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28317 \$153 \$13213 \$11987 \$13367 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$28318 \$153 \$13129 \$12353 \$12982 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28320 \$153 \$13045 \$13063 \$12093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28323 \$153 \$12987 \$13063 \$12003 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28324 \$16 \$12095 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28325 \$16 \$12093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28326 \$16 \$11987 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28327 \$153 \$13130 \$11949 \$13113 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$28328 \$16 \$12003 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28330 \$153 \$13114 \$12842 \$12093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28332 \$16 \$11949 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28334 \$16 \$12158 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28335 \$153 \$13114 \$12229 \$12924 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28336 \$16 \$12093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28337 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$28338 \$153 \$13191 \$12842 \$12230 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28339 \$153 \$13064 \$12842 \$12095 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28341 \$16 \$12230 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28342 \$153 \$13064 \$12353 \$12924 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28343 \$16 \$12095 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28344 \$16 \$12093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28345 \$153 \$13250 \$11888 \$13192 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$28346 \$153 \$13046 \$12874 \$12236 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28347 \$153 \$13115 \$12013 \$13184 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$28350 \$153 \$12844 \$12874 \$12230 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28351 \$16 \$11721 \$12779 \$13184 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$28352 \$153 \$13193 \$13115 \$12093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28353 \$153 \$13131 \$13115 \$12003 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28356 \$16 \$11721 \$16 \$153 \$13194 VNB sky130_fd_sc_hd__inv_1
X$28357 \$153 \$13157 \$12720 \$12236 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28358 \$153 \$12990 \$12720 \$12152 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28359 \$16 \$12294 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28360 \$153 \$13195 \$13188 \$12093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28361 \$16 \$12152 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28362 \$16 \$12236 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28363 \$16 \$11721 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28365 \$16 \$11800 \$12897 \$13104 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$28366 \$153 \$13188 \$11897 \$13104 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$28367 \$153 \$13185 \$13188 \$12003 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28369 \$153 \$13132 \$12875 \$12294 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28370 \$16 \$11800 \$16 \$153 \$13216 VNB sky130_fd_sc_hd__inv_1
X$28371 \$16 \$12003 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28373 \$16 \$11800 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28375 \$153 \$13132 \$12208 \$12926 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28376 \$16 \$12294 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28378 \$153 \$13066 \$12875 \$12152 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28379 \$153 \$13116 \$12875 \$12230 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28381 \$153 \$13066 \$12209 \$12926 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28382 \$16 \$12152 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28383 \$16 \$12230 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28384 \$16 \$11637 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28386 \$153 \$13158 \$12921 \$12158 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28388 \$153 \$13133 \$12921 \$12093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28389 \$16 \$12158 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28390 \$153 \$13116 \$12412 \$12926 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28393 \$16 \$12093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28394 \$16 \$12093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28395 \$16 \$11814 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28398 \$153 \$13047 \$12921 \$12095 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28399 \$153 \$13186 \$12921 \$12230 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28400 \$16 \$12230 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28401 \$16 \$12095 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28402 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$28403 \$16 \$11267 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28405 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$28406 \$16 \$12158 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28407 \$16 \$10974 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28408 \$153 \$13159 \$12993 \$12158 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28409 \$153 \$13134 \$12993 \$12152 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28410 \$153 \$13134 \$12209 \$13108 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28412 \$153 \$13068 \$12208 \$13108 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28415 \$16 \$12093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28417 \$153 \$13135 \$12993 \$12095 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28418 \$153 \$13160 \$12993 \$12093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28419 \$16 \$12095 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28420 \$153 \$13135 \$12353 \$13108 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28422 \$16 \$11289 \$12922 \$13117 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$28424 \$153 \$13187 \$12134 \$13108 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28425 \$153 \$13118 \$11432 \$13117 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$28427 \$153 \$13161 \$13118 \$12044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28429 \$153 \$13069 \$13118 \$12295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28430 \$16 \$12044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28432 \$153 \$13161 \$12068 \$13105 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28433 \$153 \$13069 \$12155 \$13105 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28434 \$16 \$11289 \$16 \$153 \$13105 VNB sky130_fd_sc_hd__inv_1
X$28435 \$153 \$13136 \$13118 \$12241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28436 \$16 \$11289 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28438 \$153 \$13162 \$13118 \$12083 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28440 \$153 \$13070 \$12877 \$12241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28441 \$153 \$13162 \$12174 \$13105 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28442 \$153 \$13136 \$12363 \$13105 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28443 \$153 \$13070 \$12363 \$12928 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28444 \$16 \$11757 \$12922 \$13221 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$28445 \$153 \$13137 \$12848 \$12295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28446 \$16 \$11757 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28448 \$16 \$11757 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28450 \$16 \$11721 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28451 \$153 \$13196 \$12174 \$13222 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28452 \$153 \$13137 \$12155 \$12781 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28453 \$153 \$13119 \$12848 \$12259 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28454 \$16 \$12295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28455 \$16 \$11274 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28456 \$16 \$11794 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28459 \$153 \$13119 \$12307 \$12781 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28460 \$16 \$11721 \$12922 \$13189 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$28461 \$16 \$12259 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28462 \$153 \$13138 \$12997 \$12296 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28463 \$153 \$13163 \$12997 \$12160 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28464 \$16 \$12044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28465 \$16 \$12296 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28468 \$153 \$13106 \$12997 \$12101 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28469 \$153 \$13138 \$12359 \$13071 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28470 \$16 \$12160 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28471 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$28472 \$153 \$13106 \$12476 \$13071 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28473 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$28474 \$16 \$12101 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28475 \$153 \$13164 \$12997 \$12044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28477 \$153 \$13073 \$12997 \$12259 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28479 \$153 \$13164 \$12068 \$13071 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28480 \$153 \$13073 \$12307 \$13071 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28481 \$16 \$12259 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28482 \$153 \$13072 \$12155 \$13071 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28483 \$16 \$12044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28485 \$153 \$13190 \$11637 \$13197 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$28487 \$153 \$13042 \$11897 \$13074 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$28488 \$16 \$11637 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28490 \$153 \$13165 \$13190 \$12101 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28491 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$28493 \$16 \$12101 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28495 \$153 \$13036 \$13042 \$12259 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28496 \$16 \$11800 \$16 \$153 \$13049 VNB sky130_fd_sc_hd__inv_1
X$28498 \$153 \$13166 \$13042 \$12295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28499 \$16 \$12259 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28500 \$153 \$13139 \$13042 \$12160 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28501 \$16 \$12295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28505 \$153 \$13139 \$12028 \$13049 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28507 \$153 \$13140 \$13042 \$12296 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28508 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$28510 \$153 \$13167 \$13042 \$12083 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28511 \$16 \$12296 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28513 \$16 \$12241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28515 \$153 \$13141 \$13042 \$12241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28516 \$153 \$13140 \$12359 \$13049 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28517 \$153 \$13167 \$12174 \$13049 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28518 \$153 \$13142 \$12956 \$12083 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28519 \$16 \$12083 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28521 \$16 \$12296 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28525 \$153 \$13142 \$12174 \$13051 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28526 \$153 \$13050 \$12956 \$12101 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28528 \$153 \$13168 \$12999 \$12259 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28529 \$16 \$12083 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28530 \$16 \$12101 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28531 \$16 \$11267 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28532 \$16 \$12083 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28534 \$153 \$13076 \$12028 \$13077 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28535 \$153 \$13168 \$12307 \$13077 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28536 \$16 \$12259 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28538 \$153 \$13078 \$12999 \$12083 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28539 \$16 \$12296 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28540 \$153 \$13169 \$12999 \$12044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28541 \$16 \$12083 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28543 \$153 \$13078 \$12174 \$13077 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28544 \$16 \$12044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28545 \$16 \$12241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28546 \$153 \$13169 \$12068 \$13077 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28547 \$153 \$13079 \$12068 \$12881 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28548 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$28551 \$153 \$12882 \$12264 \$12690 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28552 \$16 \$12164 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28553 \$153 \$13170 \$12984 \$12164 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28555 \$153 \$13080 \$12984 \$12297 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28557 \$153 \$13170 \$12217 \$12932 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28558 \$153 \$13080 \$12582 \$12932 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28559 \$153 \$13198 \$12309 \$12932 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28560 \$153 \$13081 \$12984 \$12219 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28564 \$153 \$13199 \$12984 \$12298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28565 \$153 \$13081 \$12110 \$12932 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28566 \$16 \$12298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28567 \$16 \$11451 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28568 \$16 \$11399 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28569 \$153 \$13226 \$12110 \$13200 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28570 \$16 \$11578 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28571 \$16 \$12233 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28573 \$153 \$13082 \$12985 \$12233 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28575 \$153 \$13171 \$12985 \$12219 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28576 \$153 \$13082 \$12603 \$12935 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28577 \$153 \$13171 \$12110 \$12935 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28579 \$16 \$12164 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28581 \$153 \$13005 \$12985 \$12164 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28582 \$153 \$13201 \$12985 \$12297 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28583 \$153 \$13083 \$12234 \$12935 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28584 \$16 \$12297 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28585 \$153 \$13258 \$11842 \$13143 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$28587 \$16 \$12571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28589 \$16 \$11930 \$12634 \$13143 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$28590 \$16 \$12297 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28592 \$153 \$13172 \$12856 \$12571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28593 \$153 \$13084 \$12856 \$12297 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28594 \$16 \$12032 \$12634 \$13202 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$28595 \$16 \$12115 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28596 \$16 \$11930 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28598 \$16 \$12115 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28601 \$153 \$13085 \$12856 \$12115 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28603 \$153 \$13052 \$12856 \$12298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28604 \$153 \$13085 \$12234 \$12832 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28605 \$16 \$12032 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28606 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$28607 \$16 \$12233 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28608 \$153 \$13173 \$12916 \$12233 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28609 \$16 \$12297 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28611 \$153 \$13144 \$12916 \$12297 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28612 \$153 \$13144 \$12582 \$12833 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28614 \$16 \$12219 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28615 \$153 \$13145 \$12916 \$12219 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28616 \$16 \$11945 \$12634 \$13228 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$28617 \$16 \$11945 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28619 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$28620 \$153 \$13145 \$12110 \$12833 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28621 \$153 \$13053 \$12916 \$12298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28622 \$16 \$11945 \$16 \$153 \$13203 VNB sky130_fd_sc_hd__inv_1
X$28624 \$153 \$13204 \$13054 \$12115 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28625 \$16 \$11945 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28626 \$16 \$11776 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28628 \$153 \$13054 \$11776 \$13086 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$28630 \$16 \$11627 \$16 \$153 \$12648 VNB sky130_fd_sc_hd__inv_1
X$28632 \$16 \$12571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28633 \$153 \$13230 \$12917 \$12571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28634 \$16 \$12219 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28635 \$153 \$13147 \$12917 \$12219 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28637 \$16 \$12219 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28639 \$153 \$13146 \$12917 \$12297 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28640 \$153 \$13147 \$12110 \$12863 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28641 \$153 \$13174 \$12917 \$12233 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28642 \$16 \$12233 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28643 \$16 \$11798 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28644 \$16 \$12820 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28645 \$16 \$12219 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28648 \$153 \$13120 \$12264 \$13109 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28649 \$16 \$12820 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28650 \$153 \$13260 \$11921 \$13088 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$28651 \$16 \$11483 \$12820 \$13089 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$28652 \$153 \$13148 \$13110 \$12219 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28653 \$153 \$13174 \$12603 \$12863 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28654 \$16 \$11483 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28656 \$153 \$13148 \$12110 \$13205 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28657 \$153 \$13110 \$11946 \$13089 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$28658 \$16 \$11483 \$16 \$153 \$13205 VNB sky130_fd_sc_hd__inv_1
X$28659 \$153 \$13176 \$13175 \$12219 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28660 \$153 \$13010 \$12264 \$12863 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28661 \$16 \$11946 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28664 \$153 \$13121 \$13175 \$12298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28665 \$16 \$12298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28666 \$153 \$13121 \$12165 \$13149 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28668 \$16 \$11747 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28669 \$153 \$13175 \$11747 \$13122 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$28670 \$153 \$13091 \$12165 \$12836 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28672 \$16 \$12115 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28674 \$153 \$13395 \$11385 \$13123 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$28675 \$153 \$13177 \$13175 \$12115 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28676 \$16 \$11546 \$12820 \$13123 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$28677 \$153 \$13177 \$12234 \$13149 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28678 \$16 \$11459 \$16 \$153 \$13149 VNB sky130_fd_sc_hd__inv_1
X$28679 \$16 \$12820 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28682 \$16 \$11983 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28683 \$16 \$12287 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28686 \$16 \$12299 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28687 \$153 \$13150 \$13012 \$11983 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28688 \$153 \$13178 \$13012 \$12299 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28689 \$16 \$11546 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28690 \$153 \$13178 \$12371 \$13093 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28692 \$153 \$13092 \$11942 \$13093 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28695 \$153 \$13179 \$13012 \$12120 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28696 \$153 \$13150 \$11881 \$13093 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28697 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$28698 \$16 \$12162 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28699 \$153 \$12970 \$12182 \$12650 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28700 \$153 \$13179 \$12182 \$13093 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28701 \$16 \$12120 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28702 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$28704 \$16 \$11983 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28705 \$153 \$13151 \$13094 \$12120 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28706 \$153 \$13055 \$13094 \$11983 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28708 \$153 \$13152 \$11842 \$13124 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$28709 \$153 \$13151 \$12182 \$13056 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28712 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$28713 \$16 \$12120 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28714 \$16 \$12009 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28715 \$153 \$13153 \$13152 \$12120 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28716 \$153 \$13180 \$12009 \$13125 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$28717 \$153 \$13153 \$12182 \$13058 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28718 \$16 \$11772 \$12747 \$13125 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$28719 \$16 \$11772 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28721 \$16 \$11930 \$16 \$153 \$13058 VNB sky130_fd_sc_hd__inv_1
X$28722 \$16 \$11930 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28724 \$16 \$12299 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28726 \$16 \$11772 \$16 \$153 \$13181 VNB sky130_fd_sc_hd__inv_1
X$28727 \$153 \$13095 \$12227 \$12838 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28728 \$153 \$13040 \$12119 \$12838 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28729 \$153 \$13154 \$12888 \$12299 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28730 \$153 \$13206 \$11881 \$13181 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28732 \$16 \$12287 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28734 \$153 \$13154 \$12371 \$12838 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28735 \$153 \$13059 \$12888 \$12287 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28736 \$153 \$13015 \$12889 \$12351 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28738 \$153 \$13096 \$12182 \$12825 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28739 \$16 \$11945 \$12747 \$13207 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$28741 \$16 \$12032 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28742 \$16 \$12303 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28743 \$16 \$12299 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28744 \$153 \$13060 \$12889 \$12303 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28745 \$153 \$13097 \$12889 \$12299 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28746 \$16 \$12169 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28747 \$153 \$13097 \$12371 \$12825 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28748 \$16 \$11945 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28749 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$28751 \$16 \$12303 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28752 \$16 \$12299 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28753 \$153 \$13098 \$12890 \$12299 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28754 \$153 \$13061 \$12890 \$12303 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28756 \$153 \$13098 \$12371 \$12907 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28757 \$16 \$12287 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28758 \$153 \$13099 \$12890 \$12287 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28760 \$153 \$13100 \$12890 \$12120 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28761 \$16 \$12351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28762 \$16 \$11983 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28763 \$153 \$13126 \$11747 \$12976 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$28764 \$153 \$13100 \$12182 \$12907 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28765 \$16 \$12303 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28769 \$153 \$13155 \$13126 \$11983 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28770 \$153 \$13182 \$13126 \$12384 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28771 \$153 \$13101 \$12119 \$12750 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28772 \$153 \$13208 \$12182 \$13209 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28774 \$16 \$12384 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28775 \$16 \$11459 \$16 \$153 \$13209 VNB sky130_fd_sc_hd__inv_1
X$28777 \$16 \$11483 \$12678 \$13127 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$28778 \$153 \$13210 \$13156 \$12384 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28779 \$153 \$13156 \$11921 \$12979 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$28780 \$153 \$13155 \$11881 \$13209 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28782 \$153 \$13265 \$11946 \$13127 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$28783 \$16 \$11946 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28786 \$16 \$11983 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28787 \$153 \$13128 \$13020 \$11983 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28788 \$16 \$11172 \$16 \$153 \$13107 VNB sky130_fd_sc_hd__inv_1
X$28789 \$153 \$13128 \$11881 \$13107 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28790 \$153 \$13102 \$12182 \$13107 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28791 \$153 \$13062 \$13020 \$12287 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28794 \$153 \$13103 \$11942 \$13107 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28795 \$16 \$12287 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28796 \$16 \$12299 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28798 \$153 \$13111 \$13020 \$12299 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28799 \$16 \$12384 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28800 \$153 \$13183 \$13020 \$12384 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28801 \$16 \$12351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28803 \$153 \$13111 \$12371 \$13107 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28805 \$153 \$13211 \$12227 \$13107 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28806 \$153 \$11557 \$10466 \$12782 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28807 \$153 \$13183 \$12179 \$13107 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28809 \$153 \$11463 \$10815 \$12782 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28810 \$153 \$13024 \$12179 \$12980 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28812 \$16 \$12782 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28813 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$28814 \$16 \$12782 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28816 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$28817 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$28818 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$28819 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$28820 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$28821 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$28824 \$153 \$3445 \$3708 \$3766 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28825 \$153 \$3391 \$3708 \$3709 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28826 \$16 \$3709 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28827 \$16 \$3616 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28828 \$153 \$3776 \$3389 \$3765 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28829 \$16 \$3766 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28832 \$153 \$3390 \$3708 \$3616 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28833 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$28834 \$153 \$3628 \$3708 \$3473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28835 \$153 \$3286 \$3708 \$3615 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28836 \$16 \$3473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28839 \$153 \$3494 \$5151 \$3734 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$28840 \$16 \$3615 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28841 \$16 \$5151 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28842 \$153 \$3268 \$3708 \$3571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28844 \$153 \$3723 \$3495 \$3766 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28845 \$16 \$3638 \$16 \$153 \$3208 VNB sky130_fd_sc_hd__inv_1
X$28848 \$16 \$3638 \$3686 \$3900 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$28849 \$16 \$3616 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28850 \$16 \$3766 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28852 \$153 \$3844 \$3864 \$3615 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28853 \$153 \$3495 \$3767 \$3777 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$28854 \$16 \$3841 \$3686 \$3777 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$28856 \$153 \$3844 \$3307 \$3934 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28857 \$16 \$3686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28859 \$16 \$3767 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28860 \$16 \$3841 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28861 \$153 \$3735 \$3606 \$3331 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28863 \$153 \$3798 \$3497 \$3709 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28864 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$28865 \$153 \$3873 \$3394 \$3872 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28867 \$16 \$3778 \$3686 \$3768 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$28868 \$153 \$3497 \$4079 \$3768 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$28870 \$153 \$3655 \$3389 \$3426 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28871 \$16 \$3778 \$16 \$153 \$3426 VNB sky130_fd_sc_hd__inv_1
X$28872 \$153 \$3736 \$3307 \$3426 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28873 \$153 \$3836 \$3845 \$3571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28874 \$16 \$4079 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28875 \$16 \$3778 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28878 \$153 \$3873 \$3845 \$3385 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28879 \$16 \$3571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28880 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$28881 \$153 \$3737 \$3606 \$3578 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28882 \$16 \$3709 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28883 \$16 \$3385 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28885 \$16 \$3761 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28887 \$153 \$3407 \$5183 \$3738 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$28888 \$153 \$3874 \$3389 \$3872 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28890 \$153 \$3874 \$3845 \$3616 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28891 \$16 \$5183 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28892 \$16 \$3761 \$3686 \$3799 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$28893 \$153 \$3800 \$3408 \$3616 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28894 \$153 \$3408 \$5095 \$3799 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$28897 \$153 \$3801 \$3408 \$3709 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28898 \$153 \$3800 \$3389 \$3476 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28899 \$16 \$3709 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28900 \$153 \$3801 \$3606 \$3476 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28901 \$153 \$3802 \$3499 \$3616 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28902 \$16 \$3761 \$16 \$153 \$3476 VNB sky130_fd_sc_hd__inv_1
X$28903 \$16 \$3571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28906 \$153 \$3903 \$3422 \$3875 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28907 \$16 \$3616 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28909 \$153 \$3769 \$3606 \$3409 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28911 \$153 \$3846 \$3838 \$3571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28912 \$153 \$3802 \$3389 \$3409 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28913 \$16 \$3385 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28914 \$153 \$3904 \$3838 \$3615 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28916 \$16 \$3571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28918 \$153 \$3803 \$3410 \$3709 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28919 \$16 \$3615 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28920 \$16 \$3615 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28921 \$153 \$3803 \$3606 \$3334 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28922 \$16 \$3766 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28923 \$16 \$3709 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28925 \$153 \$3724 \$3410 \$3616 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28928 \$153 \$3905 \$4077 \$3615 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28929 \$153 \$3632 \$3725 \$3385 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28930 \$153 \$3847 \$3725 \$3473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28932 \$16 \$3616 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28933 \$16 \$3385 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28934 \$153 \$3739 \$3422 \$3607 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28935 \$153 \$3847 \$3540 \$3607 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28936 \$153 \$3174 \$1792 \$2634 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28937 \$16 \$3473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28939 \$153 \$3740 \$3490 \$3607 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28940 \$16 \$3906 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28941 \$16 \$3907 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28942 \$153 \$3804 \$3725 \$3766 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28943 \$16 \$3907 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28945 \$16 \$2743 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28946 \$153 \$3741 \$3389 \$3607 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28947 \$16 \$3709 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28948 \$153 \$3804 \$3478 \$3607 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28949 \$16 \$1325 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28950 \$16 \$1325 \$16 \$153 \$2576 VNB sky130_fd_sc_hd__clkbuf_2
X$28951 \$16 \$2634 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28952 \$16 \$3616 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28953 \$153 \$3591 \$3909 \$3397 \$3865 \$3866 \$3867 \$3592 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$28954 \$16 \$3766 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28955 \$16 \$1943 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28957 \$153 \$3591 \$3805 \$3448 \$3779 \$3780 \$3781 \$3592 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$28958 \$16 \$3712 \$3911 \$3742 \$204 \$16 \$153 VNB sky130_fd_sc_hd__mux2_1
X$28959 \$153 \$3591 \$3743 \$3289 \$3839 \$3811 \$3636 \$3592 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$28961 \$16 \$3310 \$16 \$153 \$3591 VNB sky130_fd_sc_hd__clkbuf_2
X$28963 \$16 \$3310 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28964 \$16 \$3241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28965 \$16 \$3783 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28966 \$16 \$3638 \$3783 \$3782 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$28967 \$153 \$3848 \$3785 \$3621 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28968 \$153 \$3412 \$3660 \$3782 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$28969 \$153 \$3848 \$3608 \$3868 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28971 \$16 \$3621 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28972 \$16 \$3783 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28973 \$16 \$3692 \$3783 \$3784 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$28974 \$153 \$3876 \$3079 \$3868 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28975 \$153 \$3713 \$5151 \$3784 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$28976 \$16 \$5151 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28977 \$153 \$3661 \$3645 \$3336 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28979 \$153 \$3806 \$3785 \$3492 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28981 \$153 \$3849 \$3785 \$3386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28983 \$153 \$3806 \$3354 \$3868 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28984 \$153 \$3849 \$3435 \$3868 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28985 \$16 \$3621 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28986 \$16 \$3386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28987 \$16 \$3492 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28988 \$153 \$3877 \$3354 \$4022 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28990 \$153 \$3662 \$3713 \$3543 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$28992 \$16 \$3767 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28993 \$153 \$3878 \$3435 \$4068 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$28994 \$153 \$3502 \$3767 \$3840 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$28995 \$16 \$3841 \$3783 \$3840 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$28996 \$16 \$3543 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28997 \$16 \$3783 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$28999 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$29000 \$16 \$3543 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29001 \$16 \$3841 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29002 \$153 \$3771 \$3502 \$3543 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29003 \$153 \$3771 \$3556 \$3337 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29004 \$153 \$3644 \$3502 \$3620 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29005 \$16 \$3761 \$3783 \$3912 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$29006 \$16 \$3841 \$16 \$153 \$3337 VNB sky130_fd_sc_hd__inv_1
X$29008 \$153 \$3807 \$3413 \$3543 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29009 \$16 \$3620 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29010 \$16 \$3783 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29011 \$16 \$3761 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29012 \$16 \$3879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29013 \$153 \$3850 \$3955 \$3573 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29014 \$153 \$3808 \$3413 \$3620 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29015 \$16 \$3573 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29018 \$153 \$3808 \$3645 \$3339 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29019 \$16 \$3761 \$16 \$153 \$3339 VNB sky130_fd_sc_hd__inv_1
X$29020 \$16 \$3714 \$3783 \$3786 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$29021 \$153 \$3807 \$3556 \$3339 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29022 \$153 \$3542 \$5183 \$3786 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$29023 \$16 \$3783 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29025 \$153 \$3880 \$3079 \$3881 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29026 \$16 \$3761 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29029 \$153 \$3698 \$3608 \$3506 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29030 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$29031 \$16 \$3842 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29032 \$153 \$3851 \$3869 \$3492 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29033 \$16 \$3714 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29034 \$153 \$3727 \$3542 \$3620 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29035 \$16 \$3492 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29036 \$16 \$4107 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29038 \$153 \$3744 \$3101 \$3506 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29039 \$153 \$3882 \$3435 \$3881 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29040 \$16 \$3620 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29041 \$153 \$3851 \$3354 \$3881 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29042 \$153 \$3809 \$3493 \$3620 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29044 \$16 \$3997 \$16 \$153 \$3340 VNB sky130_fd_sc_hd__inv_1
X$29045 \$153 \$3883 \$3435 \$3884 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29047 \$153 \$3810 \$3493 \$3543 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29048 \$153 \$3809 \$3645 \$3340 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29049 \$16 \$3949 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29050 \$153 \$3574 \$3949 \$3885 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$29051 \$16 \$3620 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29052 \$153 \$3745 \$3608 \$3340 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29053 \$16 \$3543 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29055 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$29056 \$16 \$3886 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29057 \$16 \$3658 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29058 \$153 \$3887 \$3079 \$3884 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29059 \$153 \$3728 \$3574 \$3620 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29060 \$153 \$3648 \$3574 \$3621 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29061 \$16 \$3658 \$16 \$153 \$3436 VNB sky130_fd_sc_hd__inv_1
X$29062 \$16 \$3620 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29063 \$16 \$3658 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29065 \$16 \$3573 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29066 \$16 \$3621 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29067 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$29068 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$29070 \$153 \$3812 \$3787 \$3492 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29071 \$153 \$3729 \$3787 \$3573 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29072 \$16 \$3492 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29073 \$16 \$3572 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29074 \$16 \$3772 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29075 \$16 \$3573 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29077 \$16 \$3939 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29079 \$16 \$3480 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29080 \$16 \$3907 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29081 \$153 \$3813 \$3787 \$3620 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29082 \$16 \$3907 \$16 \$153 \$3585 VNB sky130_fd_sc_hd__inv_1
X$29083 \$153 \$3888 \$3787 \$3480 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29084 \$153 \$3813 \$3645 \$3585 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29085 \$16 \$3620 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29086 \$16 \$3645 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29087 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29088 \$153 \$3711 \$1482 \$3919 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29090 \$153 \$1367 \$3386 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$29091 \$153 \$3888 \$3504 \$3585 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29092 \$153 \$3811 \$1482 \$3939 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29093 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29094 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29096 \$153 \$3276 \$3852 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$29097 \$153 \$3244 \$3814 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$29098 \$16 \$3276 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29099 \$16 \$3272 \$3916 \$3128 \$721 \$16 \$153 VNB sky130_fd_sc_hd__mux2_1
X$29101 \$16 \$1367 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29103 \$153 \$3789 \$3788 \$3762 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29104 \$153 \$3333 \$3791 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$29105 \$153 \$3288 \$3792 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$29106 \$16 \$3288 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29107 \$16 \$2092 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29110 \$16 \$1868 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29111 \$153 \$3853 \$3958 \$3852 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29112 \$16 \$2026 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29113 \$16 \$1993 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29115 \$16 \$1879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29116 \$153 \$3917 \$3919 \$3762 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29117 \$153 \$3853 \$3763 \$3762 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29118 \$16 \$1665 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29119 \$16 \$1712 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29120 \$16 \$3792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29121 \$16 \$3852 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29123 \$153 \$3699 \$3715 \$3792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29124 \$153 \$3815 \$3715 \$3852 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29126 \$153 \$3815 \$3763 \$3160 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29128 \$16 \$3814 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29129 \$153 \$3293 \$3715 \$3814 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29130 \$16 \$3357 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29133 \$16 \$3889 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29135 \$16 \$3852 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29136 \$153 \$3746 \$3788 \$3890 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29137 \$16 \$3731 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29138 \$16 \$3814 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29139 \$153 \$3816 \$3790 \$3814 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29140 \$153 \$3854 \$3790 \$3852 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29143 \$16 \$3791 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29144 \$153 \$3854 \$3763 \$3890 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29145 \$153 \$3817 \$3790 \$3791 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29146 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$29148 \$16 \$3731 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29149 \$153 \$3818 \$3622 \$3731 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29151 \$153 \$3818 \$3788 \$3732 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29153 \$16 \$3791 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29154 \$153 \$3855 \$3622 \$3791 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29155 \$153 \$3819 \$3622 \$3792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29156 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$29157 \$153 \$3855 \$3919 \$3732 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29158 \$16 \$3792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29159 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$29162 \$16 \$3731 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29163 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$29164 \$153 \$3562 \$1712 \$3162 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29166 \$16 \$3792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29167 \$153 \$3856 \$3717 \$3792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29168 \$153 \$3820 \$3717 \$3731 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29169 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$29171 \$153 \$3747 \$3651 \$3773 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29172 \$153 \$3856 \$3939 \$3773 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29173 \$153 \$3748 \$3763 \$3773 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29175 \$153 \$3857 \$3670 \$3792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29176 \$153 \$3820 \$3788 \$3773 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29178 \$16 \$3792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29180 \$153 \$3821 \$3670 \$3814 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29181 \$16 \$3814 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29182 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$29183 \$153 \$3821 \$3651 \$3891 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29184 \$153 \$3671 \$3788 \$3891 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29185 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$29186 \$16 \$3814 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29187 \$153 \$3650 \$3649 \$3814 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29188 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$29190 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$29191 \$16 \$3792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29192 \$153 \$3923 \$3858 \$3609 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29193 \$153 \$3750 \$3763 \$3609 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29194 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$29195 \$153 \$3672 \$3788 \$3609 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29196 \$16 \$3792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29197 \$16 \$3889 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29198 \$153 \$3733 \$3718 \$3889 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29201 \$153 \$3774 \$3718 \$3792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29202 \$16 \$3814 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29203 \$153 \$3611 \$3718 \$3814 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29204 \$153 \$3751 \$3763 \$3610 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29205 \$16 \$3418 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29208 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29209 \$153 \$3892 \$3716 \$3610 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29210 \$153 \$3653 \$1482 \$3986 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29211 \$16 \$3822 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29212 \$153 \$3859 \$3718 \$3791 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29213 \$153 \$3774 \$3939 \$3610 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29215 \$153 \$3859 \$3919 \$3610 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29218 \$153 \$3530 \$3823 \$3312 \$3822 \$3754 \$3675 \$3511 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$29219 \$153 \$3689 \$1482 \$3860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29220 \$153 \$3510 \$1482 \$3893 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29221 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29222 \$16 \$3312 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29224 \$16 \$3860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29226 \$16 \$4276 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29227 \$16 \$3893 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29228 \$153 \$3243 \$3826 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$29229 \$153 \$3793 \$3676 \$3461 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29230 \$153 \$3794 \$3986 \$3461 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29231 \$153 \$3439 \$3898 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$29233 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29234 \$16 \$3439 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29235 \$16 \$2000 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29237 \$153 \$3824 \$3795 \$3721 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29238 \$153 \$3894 \$3860 \$3586 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29239 \$16 \$3199 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29240 \$153 \$3200 \$3602 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$29242 \$16 \$3508 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29243 \$16 \$3721 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29244 \$16 \$3898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29245 \$153 \$3825 \$3795 \$3691 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29246 \$16 \$3200 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29247 \$153 \$3843 \$3719 \$3586 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29248 \$153 \$3843 \$3795 \$3680 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29250 \$153 \$3825 \$3142 \$3586 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29251 \$16 \$3826 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29252 \$153 \$3926 \$3705 \$3826 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29253 \$16 \$3680 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29255 \$153 \$3720 \$3680 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$29256 \$16 \$3870 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29259 \$16 \$3602 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29260 \$16 \$4129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29261 \$153 \$3827 \$3705 \$3602 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29262 \$153 \$3896 \$3860 \$3895 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29263 \$153 \$3794 \$3705 \$4129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29264 \$16 \$3680 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29265 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$29267 \$16 \$3602 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29268 \$153 \$3756 \$3142 \$3775 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29269 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$29271 \$16 \$3721 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29272 \$153 \$3928 \$3796 \$3721 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29273 \$153 \$3828 \$3796 \$3602 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29274 \$16 \$3929 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29278 \$16 \$4057 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29279 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$29280 \$153 \$3829 \$3796 \$4057 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29282 \$153 \$3897 \$4414 \$3612 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29283 \$153 \$3861 \$3860 \$3612 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29285 \$153 \$3757 \$3676 \$3612 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29286 \$153 \$3830 \$3142 \$3612 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29289 \$16 \$3691 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29290 \$153 \$3830 \$3623 \$3691 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29291 \$153 \$3861 \$3623 \$3898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29292 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$29293 \$16 \$3898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29294 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$29295 \$153 \$3468 \$1936 \$2931 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29297 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$29298 \$153 \$3831 \$3624 \$3721 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29299 \$16 \$3898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29300 \$16 \$3680 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29301 \$153 \$3931 \$3624 \$3680 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29303 \$16 \$4057 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29304 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$29305 \$153 \$3831 \$3676 \$3930 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29306 \$16 \$3680 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29308 \$153 \$3758 \$4414 \$3764 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29310 \$16 \$4057 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29311 \$16 \$3721 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29312 \$153 \$3832 \$3722 \$3680 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29313 \$153 \$3833 \$3722 \$3721 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29314 \$153 \$3833 \$3676 \$3764 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29315 \$16 \$4129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29317 \$153 \$3797 \$3722 \$4129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29319 \$16 \$5002 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29320 \$16 \$3834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29322 \$153 \$3797 \$3986 \$3764 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29323 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$29324 \$16 \$4092 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29325 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$29326 \$16 \$3680 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29327 \$153 \$3862 \$3871 \$3680 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29328 \$16 \$4129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29330 \$153 \$3835 \$3625 \$4129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29331 \$153 \$3862 \$3719 \$3899 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29333 \$16 \$3834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29334 \$153 \$3382 \$2056 \$3328 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29335 \$16 \$3834 \$16 \$153 \$4171 VNB sky130_fd_sc_hd__inv_1
X$29337 \$16 \$3826 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29338 \$16 \$4057 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29341 \$16 \$3826 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29342 \$153 \$3863 \$3871 \$4057 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29343 \$153 \$4157 \$3625 \$3826 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29344 \$153 \$4380 \$3625 \$4057 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29345 \$153 \$3538 \$2269 \$3328 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29347 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$29348 \$16 \$4057 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29349 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$29350 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$29351 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$29352 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$29353 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$29354 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$29357 \$153 \$4174 \$3942 \$3709 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29358 \$153 \$3943 \$3942 \$3474 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29359 \$16 \$3709 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29361 \$153 \$4075 \$3389 \$4066 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29362 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$29364 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$29365 \$153 \$4175 \$3942 \$3385 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29366 \$153 \$4028 \$3478 \$3765 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29367 \$153 \$4174 \$3606 \$3765 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29368 \$153 \$4210 \$3394 \$4066 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29369 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$29370 \$16 \$4162 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29372 \$153 \$4100 \$3942 \$3615 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29373 \$16 \$4162 \$16 \$153 \$3765 VNB sky130_fd_sc_hd__inv_1
X$29374 \$153 \$3942 \$4083 \$4099 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$29375 \$16 \$4162 \$3686 \$4099 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$29376 \$16 \$3615 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29377 \$153 \$4101 \$3307 \$4067 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29379 \$153 \$4101 \$4158 \$3615 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29381 \$153 \$4176 \$4158 \$3709 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29382 \$153 \$4417 \$3490 \$4067 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29383 \$16 \$3616 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29384 \$153 \$4076 \$3389 \$4067 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29385 \$16 \$3615 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29387 \$153 \$4142 \$3864 \$3616 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29389 \$16 \$3709 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29391 \$153 \$4102 \$3864 \$3473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29392 \$153 \$4142 \$3389 \$3934 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29393 \$153 \$4177 \$3422 \$4067 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29394 \$153 \$4103 \$3864 \$3766 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29397 \$153 \$4102 \$3540 \$3934 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29398 \$153 \$4103 \$3478 \$3934 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29399 \$16 \$4178 \$16 \$153 \$3934 VNB sky130_fd_sc_hd__inv_1
X$29400 \$16 \$4178 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29401 \$16 \$4179 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29402 \$16 \$3766 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29404 \$153 \$4180 \$4143 \$3473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29405 \$153 \$3836 \$3422 \$3872 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29408 \$153 \$4029 \$3478 \$3872 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29409 \$16 \$3473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29410 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$29411 \$153 \$3845 \$5201 \$4104 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$29412 \$16 \$3766 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29414 \$153 \$4018 \$3845 \$3473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29416 \$16 \$3879 \$16 \$153 \$3872 VNB sky130_fd_sc_hd__inv_1
X$29418 \$16 \$5201 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29419 \$16 \$3879 \$3686 \$4104 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$29420 \$16 \$3879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29421 \$16 \$3879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29422 \$16 \$3686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29423 \$16 \$3473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29425 \$153 \$4159 \$3422 \$4328 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29426 \$153 \$4105 \$3947 \$3616 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29427 \$16 \$3766 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29428 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$29429 \$153 \$4031 \$3490 \$3875 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29430 \$16 \$3616 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29432 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$29433 \$16 \$1433 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29434 \$153 \$4105 \$3389 \$3875 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29435 \$16 \$4106 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29436 \$153 \$4032 \$3947 \$3615 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29437 \$16 \$4106 \$16 \$153 \$3875 VNB sky130_fd_sc_hd__inv_1
X$29438 \$16 \$3385 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29440 \$16 \$1433 \$16 \$153 \$4181 VNB sky130_fd_sc_hd__clkbuf_2
X$29441 \$16 \$3997 \$4144 \$4145 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$29442 \$153 \$4032 \$3307 \$3875 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29444 \$153 \$3499 \$4107 \$4145 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$29445 \$16 \$3615 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29446 \$16 \$4106 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29447 \$16 \$4107 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29448 \$153 \$4034 \$3838 \$3474 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29449 \$16 \$4146 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29450 \$16 \$3474 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29451 \$153 \$3302 \$2064 \$2743 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29454 \$153 \$4213 \$3389 \$3935 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29455 \$153 \$4034 \$3490 \$3935 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29457 \$153 \$4182 \$3478 \$3935 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29458 \$153 \$4033 \$3394 \$3935 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29459 \$16 \$3709 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29460 \$153 \$4147 \$3540 \$3935 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29461 \$153 \$4108 \$4077 \$3473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29465 \$16 \$3571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29466 \$153 \$4108 \$3540 \$4019 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29468 \$153 \$3905 \$3307 \$4019 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29469 \$153 \$4183 \$4077 \$3474 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29470 \$153 \$3173 \$2064 \$2634 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29473 \$153 \$4036 \$3478 \$4019 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29474 \$153 \$4133 \$4077 \$3616 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29475 \$16 \$3886 \$4012 \$4109 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$29476 \$16 \$3766 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29477 \$153 \$4183 \$3490 \$4019 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29478 \$153 \$3951 \$3725 \$3615 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29479 \$16 \$3616 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29482 \$153 \$153 \$3307 \$4020 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29483 \$153 \$153 \$3389 \$4020 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29484 \$153 \$153 \$3540 \$4020 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29485 \$153 \$153 \$3490 \$4020 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29486 \$153 \$153 \$3478 \$4020 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29487 \$16 \$1918 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29488 \$16 \$3780 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29489 \$16 \$4079 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29492 \$16 \$4134 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29493 \$16 \$4078 \$16 \$153 \$4110 VNB sky130_fd_sc_hd__clkbuf_2
X$29494 \$16 \$4184 \$16 \$153 \$4160 VNB sky130_fd_sc_hd__clkbuf_2
X$29495 \$16 \$4080 \$16 \$153 \$3692 VNB sky130_fd_sc_hd__clkbuf_2
X$29496 \$153 \$4081 \$4160 \$4148 \$4110 \$4215 \$16 \$16 VNB
+ sky130_fd_sc_hd__nor4b_2
X$29498 \$16 \$4081 \$16 \$153 \$3714 VNB sky130_fd_sc_hd__clkbuf_2
X$29499 \$16 \$4082 \$16 \$153 \$3761 VNB sky130_fd_sc_hd__clkbuf_2
X$29500 \$153 \$3785 \$4079 \$4038 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$29501 \$153 \$4148 \$4110 \$4161 \$4160 \$4215 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$29504 \$16 \$4162 \$3783 \$4135 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$29505 \$153 \$4111 \$4083 \$4135 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$29506 \$16 \$3783 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29508 \$153 \$4084 \$4111 \$3621 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29509 \$16 \$4083 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29510 \$153 \$4084 \$3608 \$4022 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29511 \$16 \$4162 \$16 \$153 \$4022 VNB sky130_fd_sc_hd__inv_1
X$29513 \$16 \$3621 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29515 \$16 \$3573 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29516 \$153 \$4085 \$4111 \$3543 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29517 \$153 \$4021 \$4111 \$3573 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29518 \$153 \$4185 \$3101 \$4022 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29519 \$153 \$4085 \$3556 \$4022 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29520 \$16 \$3543 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29521 \$153 \$4086 \$3504 \$4022 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29523 \$16 \$3573 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29524 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$29525 \$153 \$4186 \$4111 \$3386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29526 \$153 \$4112 \$4111 \$3620 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29528 \$153 \$4112 \$3645 \$4022 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29529 \$16 \$3620 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29532 \$153 \$4186 \$3435 \$4022 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29533 \$153 \$4187 \$3954 \$3620 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29534 \$16 \$4229 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29536 \$153 \$4040 \$3954 \$3543 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29537 \$16 \$3620 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29538 \$16 \$4229 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29539 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$29540 \$153 \$4040 \$3556 \$4068 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29542 \$153 \$4187 \$3645 \$4068 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29543 \$153 \$4041 \$3354 \$4068 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29545 \$16 \$3621 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29547 \$153 \$4188 \$3955 \$3572 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29548 \$153 \$3975 \$3079 \$4068 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29551 \$16 \$4178 \$16 \$153 \$3937 VNB sky130_fd_sc_hd__inv_1
X$29552 \$153 \$4188 \$3101 \$3937 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29554 \$153 \$4042 \$3608 \$3937 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29555 \$153 \$4189 \$3955 \$3543 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29556 \$16 \$3621 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29557 \$16 \$4178 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29558 \$16 \$5201 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29559 \$16 \$3480 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29560 \$153 \$3869 \$5201 \$4013 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$29561 \$16 \$3543 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29563 \$153 \$4189 \$3556 \$3937 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29564 \$16 \$3783 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29566 \$16 \$3879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29568 \$16 \$3573 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29569 \$153 \$4113 \$3869 \$3543 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29570 \$153 \$4190 \$3869 \$3621 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29572 \$153 \$4190 \$3608 \$3881 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29573 \$16 \$3879 \$16 \$153 \$3881 VNB sky130_fd_sc_hd__inv_1
X$29574 \$16 \$1485 \$16 \$153 \$4249 VNB sky130_fd_sc_hd__clkbuf_2
X$29575 \$153 \$4114 \$3869 \$3572 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29576 \$153 \$4113 \$3556 \$3881 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29577 \$16 \$3572 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29579 \$153 \$3493 \$4107 \$4069 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$29582 \$153 \$4114 \$3101 \$3881 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29584 \$153 \$4191 \$4163 \$3621 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29585 \$16 \$3997 \$4014 \$4069 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$29586 \$16 \$3621 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29587 \$153 \$4191 \$3608 \$4164 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29589 \$153 \$4115 \$3956 \$3621 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29590 \$153 \$4192 \$4163 \$3480 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29591 \$153 \$4115 \$3608 \$3884 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29592 \$16 \$3886 \$3957 \$4193 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$29594 \$153 \$4044 \$3956 \$3620 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29596 \$153 \$4136 \$3956 \$3572 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29597 \$153 \$4044 \$3645 \$3884 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29598 \$16 \$3572 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29599 \$153 \$4137 \$4194 \$3543 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29600 \$16 \$3620 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29601 \$16 \$4070 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29604 \$153 \$4116 \$4194 \$3492 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29605 \$153 \$4138 \$4194 \$3480 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29606 \$16 \$3492 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29607 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$29608 \$16 \$3543 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29609 \$153 \$4117 \$4194 \$3573 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29610 \$16 \$3480 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29613 \$153 \$4087 \$4194 \$3386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29614 \$153 \$4087 \$3435 \$4232 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29616 \$153 \$1516 \$3573 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$29617 \$16 \$3386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29618 \$16 \$3573 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29619 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$29621 \$153 \$4117 \$3079 \$4232 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29622 \$153 \$3780 \$1482 \$3962 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29623 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29625 \$153 \$1678 \$3543 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$29626 \$16 \$1516 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29629 \$153 \$153 \$3435 \$4233 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29630 \$153 \$3491 \$3960 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$29631 \$16 \$1678 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29632 \$16 \$3491 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29633 \$16 \$3244 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29634 \$16 \$3096 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29635 \$153 \$153 \$3788 \$4071 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29636 \$16 \$1471 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29637 \$16 \$1715 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29638 \$153 \$4118 \$3958 \$3792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29640 \$153 \$153 \$3962 \$4071 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29641 \$16 \$3983 \$16 \$153 \$4071 VNB sky130_fd_sc_hd__clkbuf_2
X$29642 \$153 \$4045 \$3958 \$4048 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29643 \$153 \$153 \$3651 \$4071 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29644 \$16 \$4093 \$4166 \$4149 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$29647 \$153 \$4045 \$3858 \$3762 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29648 \$153 \$3958 \$4276 \$4149 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$29649 \$16 \$3791 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29650 \$153 \$4046 \$3958 \$3889 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29651 \$16 \$3889 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29653 \$153 \$4195 \$4254 \$3814 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29655 \$153 \$4046 \$3962 \$3762 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29656 \$153 \$3715 \$4196 \$4119 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$29657 \$16 \$3870 \$4166 \$4119 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$29658 \$16 \$3960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29659 \$153 \$3701 \$3715 \$3960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29660 \$16 \$4196 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29661 \$16 \$3870 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29663 \$16 \$3731 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29665 \$153 \$4197 \$4165 \$3731 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29666 \$16 \$3870 \$16 \$153 \$3160 VNB sky130_fd_sc_hd__inv_1
X$29667 \$16 \$3870 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29668 \$16 \$4048 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29669 \$153 \$4120 \$3790 \$4048 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29670 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$29671 \$16 \$4139 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29672 \$153 \$4120 \$3858 \$3890 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29675 \$153 \$4121 \$3790 \$3889 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29676 \$16 \$4139 \$4166 \$4140 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$29677 \$16 \$4139 \$16 \$153 \$3890 VNB sky130_fd_sc_hd__inv_1
X$29678 \$153 \$4121 \$3962 \$3890 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29679 \$16 \$4139 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29680 \$153 \$3622 \$4047 \$4089 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$29681 \$16 \$3929 \$4166 \$4089 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$29684 \$16 \$3929 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29686 \$153 \$4198 \$3919 \$4167 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29687 \$153 \$3961 \$3622 \$3889 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29688 \$153 \$4150 \$3716 \$4167 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29690 \$153 \$4151 \$3651 \$4167 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29691 \$16 \$3929 \$16 \$153 \$3732 VNB sky130_fd_sc_hd__inv_1
X$29692 \$16 \$3929 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29695 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$29696 \$16 \$4048 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29697 \$153 \$4199 \$3717 \$4048 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29699 \$16 \$3889 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29700 \$153 \$4050 \$3717 \$3889 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29701 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$29702 \$153 \$4050 \$3962 \$3773 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29703 \$16 \$4011 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29704 \$16 \$4011 \$16 \$153 \$3773 VNB sky130_fd_sc_hd__inv_1
X$29706 \$16 \$4168 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29707 \$153 \$3717 \$4168 \$4122 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$29708 \$16 \$3889 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29709 \$16 \$4011 \$4015 \$4122 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$29711 \$153 \$4123 \$3670 \$3889 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29713 \$153 \$4090 \$3670 \$3960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29715 \$16 \$4011 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29717 \$153 \$4090 \$3716 \$3891 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29718 \$16 \$4258 \$16 \$153 \$3891 VNB sky130_fd_sc_hd__inv_1
X$29719 \$16 \$4258 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29721 \$16 \$4152 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29722 \$153 \$4123 \$3962 \$3891 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29723 \$153 \$3649 \$4152 \$4051 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$29724 \$153 \$4052 \$3649 \$3960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29726 \$153 \$4200 \$3649 \$3889 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29727 \$153 \$4005 \$3919 \$3609 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29728 \$16 \$4016 \$16 \$153 \$3609 VNB sky130_fd_sc_hd__inv_1
X$29729 \$153 \$4052 \$3716 \$3609 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29730 \$16 \$4016 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29731 \$16 \$3889 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29732 \$153 \$4201 \$4091 \$3889 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29734 \$153 \$4023 \$4091 \$3960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29735 \$153 \$4202 \$4091 \$3792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29736 \$16 \$3960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29737 \$16 \$3964 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29738 \$16 \$3834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29739 \$16 \$4048 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29740 \$153 \$3985 \$3763 \$4024 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29743 \$153 \$4204 \$4091 \$3731 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29744 \$153 \$4124 \$4091 \$4048 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29745 \$16 \$3731 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29746 \$153 \$4124 \$3858 \$4024 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29747 \$16 \$3986 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29749 \$16 \$4092 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29750 \$16 \$4125 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29752 \$16 \$4092 \$4015 \$4153 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$29753 \$16 \$4092 \$16 \$153 \$4024 VNB sky130_fd_sc_hd__inv_1
X$29754 \$153 \$4053 \$3919 \$4024 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29755 \$153 \$4091 \$4125 \$4153 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$29756 \$16 \$3814 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29757 \$153 \$153 \$3860 \$3941 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29759 \$16 \$3086 \$4203 \$3753 \$3462 \$16 \$153 VNB sky130_fd_sc_hd__mux2_1
X$29760 \$153 \$153 \$3986 \$3941 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29762 \$153 \$153 \$4414 \$3941 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29764 \$153 \$153 \$3676 \$3941 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29765 \$16 \$3086 \$4141 \$3823 \$3679 \$16 \$153 VNB sky130_fd_sc_hd__mux2_1
X$29766 \$153 \$153 \$3142 \$3941 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29768 \$16 \$3826 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29769 \$153 \$4154 \$3860 \$3461 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29770 \$16 \$4093 \$3988 \$4054 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$29772 \$153 \$4055 \$4094 \$3826 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29773 \$153 \$4205 \$4094 \$4057 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29774 \$153 \$4055 \$3893 \$4072 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29775 \$153 \$4205 \$4414 \$4072 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29776 \$16 \$4093 \$16 \$153 \$3586 VNB sky130_fd_sc_hd__inv_1
X$29779 \$153 \$4056 \$4094 \$4129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29780 \$153 \$4027 \$4094 \$3602 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29781 \$153 \$4056 \$3986 \$4072 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29782 \$16 \$3691 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29783 \$16 \$3602 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29784 \$16 \$4057 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29786 \$153 \$4017 \$4126 \$4308 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$29787 \$16 \$4129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29790 \$16 \$3870 \$3988 \$3966 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$29791 \$153 \$4059 \$4017 \$4057 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29792 \$153 \$3987 \$3986 \$3586 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29793 \$153 \$4169 \$3893 \$3895 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29794 \$16 \$4057 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29795 \$16 \$4126 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29796 \$16 \$3602 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29797 \$153 \$4060 \$4017 \$3602 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29800 \$153 \$4058 \$3676 \$3895 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29801 \$153 \$4170 \$3719 \$3895 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29802 \$153 \$4060 \$3565 \$3895 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29803 \$16 \$3929 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29804 \$16 \$4542 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29805 \$16 \$3461 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29806 \$16 \$4047 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29807 \$16 \$4129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29808 \$16 \$3826 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29809 \$153 \$4206 \$4095 \$4129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29811 \$153 \$4127 \$4095 \$3826 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29812 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$29814 \$16 \$3721 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29815 \$16 \$3602 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29816 \$153 \$3828 \$3565 \$3775 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29817 \$153 \$4128 \$4095 \$3602 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29819 \$153 \$4207 \$4095 \$3721 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29821 \$153 \$3990 \$3893 \$3775 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29822 \$16 \$4011 \$4156 \$4155 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$29823 \$153 \$4073 \$3719 \$3612 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29824 \$153 \$3623 \$4168 \$4155 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$29827 \$16 \$4129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29828 \$153 \$4130 \$3623 \$4129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29830 \$16 \$4011 \$16 \$153 \$3612 VNB sky130_fd_sc_hd__inv_1
X$29831 \$153 \$4062 \$3893 \$3612 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29832 \$153 \$3624 \$5264 \$4096 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$29833 \$16 \$4258 \$4156 \$4096 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$29834 \$16 \$5264 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29837 \$153 \$4130 \$3986 \$3612 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29838 \$16 \$4258 \$16 \$153 \$3930 VNB sky130_fd_sc_hd__inv_1
X$29839 \$153 \$3967 \$3624 \$4129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29840 \$16 \$4129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29841 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$29842 \$153 \$3991 \$3860 \$3930 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29843 \$153 \$3690 \$3142 \$3930 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29844 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$29847 \$16 \$4152 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29848 \$153 \$3722 \$4152 \$4063 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$29849 \$153 \$3931 \$3719 \$3930 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29850 \$153 \$3706 \$4414 \$3930 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29851 \$16 \$3680 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29852 \$153 \$4131 \$4268 \$3680 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29854 \$16 \$4016 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29855 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$29857 \$16 \$4125 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29858 \$153 \$4157 \$3893 \$4171 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29859 \$16 \$3898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29860 \$153 \$3871 \$4125 \$4074 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$29861 \$153 \$4064 \$3860 \$3764 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29862 \$16 \$3691 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29863 \$153 \$4208 \$4172 \$3691 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29864 \$16 \$4092 \$4156 \$4074 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$29867 \$153 \$4132 \$3871 \$3691 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29868 \$153 \$4208 \$3142 \$4173 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29869 \$16 \$3691 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29870 \$153 \$4132 \$3142 \$3899 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29871 \$153 \$4097 \$3676 \$3899 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29872 \$153 \$4097 \$3871 \$3721 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29875 \$153 \$4209 \$4172 \$3826 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29876 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$29878 \$153 \$4209 \$3893 \$4173 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29879 \$153 \$4098 \$4414 \$4173 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29881 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$29882 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$29884 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$29885 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$29886 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$29887 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$29888 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$29889 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$29890 \$153 \$1629 \$1465 \$17 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29891 \$153 \$1520 \$1465 \$504 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29893 \$153 \$1494 \$234 \$1187 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29894 \$16 \$263 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29897 \$153 \$1603 \$1465 \$58 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29898 \$153 \$1520 \$561 \$1535 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29899 \$16 \$710 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29900 \$16 \$58 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29901 \$153 \$1603 \$30 \$1535 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29902 \$153 \$1427 \$394 \$1187 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29904 \$16 \$249 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29908 \$16 \$1496 \$1168 \$1536 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$29909 \$153 \$1604 \$1465 \$184 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29910 \$153 \$1465 \$1503 \$1536 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$29911 \$153 \$1604 \$59 \$1535 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29912 \$153 \$1497 \$349 \$1535 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29913 \$16 \$184 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29914 \$16 \$395 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29916 \$16 \$1168 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29917 \$153 \$1521 \$1257 \$395 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29918 \$16 \$1503 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29919 \$153 \$1605 \$1257 \$249 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29920 \$153 \$1521 \$394 \$1106 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29921 \$153 \$1605 \$377 \$1106 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29924 \$153 \$1546 \$1547 \$1537 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29925 \$16 \$249 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29926 \$153 \$1606 \$1326 \$249 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29927 \$153 \$970 \$394 \$783 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29928 \$16 \$249 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29929 \$153 \$1606 \$377 \$1327 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29930 \$153 \$1431 \$102 \$1327 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29932 \$153 \$1451 \$349 \$1327 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29933 \$153 \$1657 \$1326 \$58 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29934 \$153 \$1548 \$59 \$1327 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29935 \$16 \$1404 \$16 \$153 \$1327 VNB sky130_fd_sc_hd__inv_1
X$29936 \$153 \$1549 \$394 \$1250 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29937 \$16 \$184 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29938 \$153 \$1630 \$1249 \$58 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29940 \$153 \$1549 \$1249 \$395 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29941 \$16 \$1328 \$1168 \$1607 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$29942 \$153 \$1249 \$1576 \$1607 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$29943 \$153 \$1550 \$59 \$1250 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29944 \$153 \$1499 \$377 \$1250 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29946 \$153 \$1631 \$1547 \$1594 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29947 \$16 \$1348 \$1168 \$1570 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$29948 \$16 \$184 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29950 \$153 \$1608 \$1258 \$184 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29951 \$153 \$1523 \$1258 \$58 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29952 \$153 \$1608 \$59 \$1191 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29954 \$153 \$1523 \$30 \$1191 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29955 \$16 \$1348 \$16 \$153 \$1191 VNB sky130_fd_sc_hd__inv_1
X$29957 \$153 \$1524 \$1330 \$58 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29959 \$153 \$1609 \$1330 \$184 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29960 \$153 \$1524 \$30 \$1454 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29962 \$16 \$184 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29963 \$153 \$1609 \$59 \$1454 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29964 \$16 \$249 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29966 \$153 \$1571 \$1330 \$17 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29967 \$153 \$1501 \$377 \$1454 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29969 \$153 \$1571 \$102 \$1454 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29970 \$16 \$17 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29972 \$16 \$1551 \$16 \$153 \$1454 VNB sky130_fd_sc_hd__inv_1
X$29973 \$16 \$323 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29974 \$16 \$1430 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29976 \$153 \$1466 \$1352 \$249 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29977 \$153 \$1481 \$1352 \$419 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29978 \$16 \$249 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29979 \$16 \$419 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29980 \$16 \$535 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29982 \$153 \$1526 \$1352 \$58 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29983 \$16 \$380 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$29986 \$153 \$1467 \$1352 \$184 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$29987 \$153 \$1526 \$30 \$1251 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$29989 \$16 \$1552 \$454 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$29991 \$16 \$1552 \$1596 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$29992 \$16 \$1552 \$531 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$29993 \$153 \$1625 \$249 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$29994 \$16 \$1552 \$1525 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$29996 \$16 \$1502 \$16 \$153 \$1331 VNB sky130_fd_sc_hd__clkbuf_2
X$29997 \$16 \$1502 \$16 \$153 \$1552 VNB sky130_fd_sc_hd__clkbuf_2
X$29998 \$153 \$1538 \$263 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$30000 \$16 \$1502 \$16 \$153 \$1626 VNB sky130_fd_sc_hd__clkbuf_2
X$30001 \$16 \$1626 \$1553 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$30002 \$16 \$1626 \$945 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$30003 \$16 \$234 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30004 \$153 \$1436 \$419 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$30006 \$16 \$1626 \$1311 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$30007 \$16 \$1626 \$1595 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$30008 \$16 \$1538 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30009 \$153 \$1610 \$17 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$30010 \$16 \$1182 \$757 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$30012 \$16 \$1354 \$16 \$153 \$1408 VNB sky130_fd_sc_hd__clkbuf_2
X$30014 \$153 \$1572 \$1482 \$561 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30015 \$153 \$1635 \$1482 \$234 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30016 \$153 \$1573 \$1482 \$394 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30017 \$16 \$1480 \$979 \$1660 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$30018 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30019 \$16 \$1610 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30020 \$16 \$561 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30024 \$153 \$1632 \$1504 \$293 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30025 \$153 \$1693 \$1504 \$187 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30026 \$16 \$1480 \$16 \$153 \$1633 VNB sky130_fd_sc_hd__inv_1
X$30027 \$16 \$187 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30028 \$153 \$1634 \$1504 \$209 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30029 \$16 \$293 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30030 \$16 \$1503 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30031 \$16 \$1496 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30033 \$16 \$280 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30034 \$153 \$1574 \$1504 \$73 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30035 \$16 \$209 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30036 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$30037 \$153 \$1574 \$215 \$1633 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30038 \$16 \$73 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30039 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$30041 \$16 \$754 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30042 \$16 \$1845 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30043 \$153 \$1575 \$1504 \$60 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30045 \$153 \$1661 \$1504 \$212 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30046 \$16 \$212 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30048 \$153 \$1262 \$1553 \$1636 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$30049 \$16 \$60 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30050 \$16 \$1553 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30053 \$153 \$1470 \$1262 \$209 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30055 \$16 \$1348 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30056 \$153 \$1484 \$1262 \$212 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30057 \$16 \$1348 \$16 \$153 \$1333 VNB sky130_fd_sc_hd__inv_1
X$30058 \$153 \$1527 \$1262 \$73 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30059 \$16 \$209 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30060 \$16 \$212 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30063 \$16 \$1686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30064 \$153 \$1334 \$1686 \$1662 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$30065 \$153 \$1527 \$215 \$1333 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30066 \$16 \$73 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30067 \$16 \$1404 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30068 \$153 \$1611 \$1334 \$209 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30070 \$16 \$323 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30071 \$16 \$1404 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30072 \$16 \$1404 \$16 \$153 \$1393 VNB sky130_fd_sc_hd__inv_1
X$30074 \$153 \$1554 \$1895 \$1922 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30075 \$153 \$1611 \$346 \$1393 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30076 \$16 \$209 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30078 \$16 \$1576 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30079 \$153 \$1637 \$347 \$1393 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30080 \$153 \$1528 \$1334 \$187 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30081 \$16 \$323 \$1292 \$1638 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$30084 \$153 \$1421 \$1576 \$1663 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$30085 \$153 \$1529 \$1334 \$293 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30086 \$153 \$1555 \$1421 \$187 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30087 \$153 \$1529 \$35 \$1393 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30090 \$153 \$1577 \$1421 \$293 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30091 \$16 \$1328 \$16 \$153 \$1335 VNB sky130_fd_sc_hd__inv_1
X$30092 \$16 \$187 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30094 \$16 \$293 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30095 \$153 \$1612 \$1421 \$209 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30096 \$153 \$1555 \$54 \$1335 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30097 \$153 \$1439 \$104 \$1335 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30100 \$153 \$1612 \$346 \$1335 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30101 \$16 \$73 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30102 \$16 \$209 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30103 \$153 \$1556 \$1472 \$60 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30105 \$16 \$209 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30106 \$153 \$1640 \$1472 \$209 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30107 \$16 \$60 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30109 \$153 \$1639 \$1471 \$1822 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30110 \$153 \$1556 \$104 \$1410 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30111 \$153 \$1640 \$346 \$1410 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30112 \$16 \$1508 \$946 \$1363 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$30114 \$153 \$1641 \$35 \$1410 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30115 \$16 \$505 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30117 \$153 \$1530 \$1472 \$73 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30119 \$153 \$1486 \$1472 \$187 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30120 \$153 \$1530 \$215 \$1410 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30121 \$16 \$187 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30123 \$153 \$1539 \$60 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$30124 \$16 \$73 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30125 \$16 \$18 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30128 \$153 \$1544 \$187 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$30129 \$16 \$1539 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30130 \$16 \$1354 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30131 \$16 \$1354 \$16 \$153 \$1487 VNB sky130_fd_sc_hd__clkbuf_2
X$30132 \$153 \$153 \$54 \$1487 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30133 \$16 \$1544 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30134 \$16 \$691 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30135 \$153 \$153 \$215 \$1487 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30137 \$153 \$153 \$346 \$1487 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30138 \$153 \$153 \$35 \$1487 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30139 \$153 \$1295 \$346 \$1411 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30140 \$153 \$1365 \$35 \$1411 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30141 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$30142 \$16 \$104 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30145 \$16 \$35 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30146 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30147 \$153 \$1578 \$1482 \$104 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30149 \$16 \$1610 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30150 \$16 \$1488 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30151 \$153 \$1610 \$273 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$30152 \$153 \$1222 \$253 \$1051 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30153 \$153 \$1579 \$1482 \$347 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30156 \$16 \$1625 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30157 \$153 \$1642 \$1613 \$1540 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30158 \$153 \$1625 \$82 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$30159 \$153 \$1557 \$1558 \$1540 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30160 \$16 \$347 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30161 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30163 \$153 \$2364 \$1482 \$559 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30164 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30165 \$16 \$346 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30167 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30168 \$153 \$1664 \$1482 \$44 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30169 \$153 \$1597 \$1482 \$112 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30170 \$16 \$44 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30172 \$16 \$424 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30173 \$153 \$1643 \$1183 \$424 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30174 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30175 \$153 \$1443 \$266 \$1252 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30176 \$153 \$1509 \$389 \$1252 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30177 \$153 \$1644 \$1613 \$1679 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30178 \$16 \$112 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30179 \$153 \$1643 \$353 \$1252 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30181 \$153 \$1559 \$388 \$1252 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30182 \$16 \$1543 \$16 \$153 \$1252 VNB sky130_fd_sc_hd__inv_1
X$30183 \$16 \$241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30184 \$153 \$1531 \$1268 \$82 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30186 \$153 \$1614 \$1268 \$241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30187 \$153 \$1511 \$389 \$1396 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30189 \$153 \$1614 \$388 \$1396 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30190 \$153 \$1531 \$44 \$1396 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30191 \$16 \$241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30193 \$153 \$1615 \$1338 \$273 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30194 \$153 \$1444 \$266 \$1396 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30195 \$16 \$273 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30198 \$16 \$1585 \$1446 \$1580 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$30199 \$153 \$1598 \$44 \$1456 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30200 \$153 \$1370 \$112 \$1541 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30201 \$153 \$1582 \$389 \$1456 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30202 \$153 \$1513 \$266 \$1541 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30203 \$153 \$1369 \$559 \$1541 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30204 \$153 \$1581 \$1253 \$273 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30207 \$153 \$1645 \$388 \$1541 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30208 \$153 \$1581 \$389 \$1541 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30209 \$16 \$273 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30210 \$153 \$1560 \$353 \$1541 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30211 \$16 \$424 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30212 \$16 \$1446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30214 \$16 \$424 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30215 \$16 \$1446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30216 \$16 \$145 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30217 \$16 \$1566 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30218 \$153 \$1646 \$1270 \$145 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30220 \$16 \$273 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30221 \$16 \$82 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30222 \$153 \$1582 \$1270 \$273 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30223 \$153 \$1299 \$21 \$1541 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30224 \$153 \$1561 \$266 \$1412 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30225 \$16 \$1518 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30226 \$16 \$1647 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30229 \$153 \$1562 \$1558 \$1542 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30230 \$16 \$145 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30231 \$153 \$1561 \$1254 \$145 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30232 \$153 \$1339 \$1254 \$82 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30233 \$153 \$1563 \$1254 \$241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30234 \$16 \$241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30237 \$16 \$1758 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30238 \$153 \$1563 \$388 \$1412 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30239 \$153 \$1648 \$353 \$1412 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30240 \$16 \$1446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30241 \$16 \$1446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30242 \$16 \$1599 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30243 \$16 \$241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30244 \$16 \$1649 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30245 \$153 \$1532 \$1320 \$241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30246 \$153 \$1583 \$44 \$1240 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30249 \$16 \$1599 \$16 \$153 \$1240 VNB sky130_fd_sc_hd__inv_1
X$30250 \$153 \$1716 \$353 \$1240 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30251 \$153 \$1583 \$1320 \$82 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30252 \$153 \$1532 \$388 \$1240 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30253 \$16 \$1475 \$1446 \$1584 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$30254 \$16 \$1599 \$1446 \$1717 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$30256 \$16 \$273 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30259 \$153 \$1533 \$1424 \$424 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30260 \$153 \$1617 \$1424 \$273 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30261 \$153 \$1617 \$389 \$1229 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30262 \$153 \$1533 \$353 \$1229 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30263 \$16 \$57 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30264 \$153 \$1515 \$44 \$1229 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30266 \$153 \$1448 \$559 \$1229 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30268 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30269 \$153 \$1650 \$1482 \$703 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30270 \$16 \$23 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30273 \$16 \$1673 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30274 \$16 \$703 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30275 \$153 \$1673 \$509 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$30276 \$16 \$1539 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30277 \$16 \$1543 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30278 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30280 \$16 \$1585 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30281 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30282 \$16 \$1543 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30284 \$16 \$902 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30285 \$153 \$1665 \$1482 \$223 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30286 \$16 \$1601 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30287 \$16 \$1544 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30288 \$153 \$1544 \$63 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$30289 \$16 \$223 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30290 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30291 \$16 \$398 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30293 \$16 \$1564 \$700 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$30295 \$16 \$1721 \$16 \$153 \$1564 VNB sky130_fd_sc_hd__clkbuf_2
X$30298 \$16 \$446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30300 \$16 \$1564 \$723 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$30301 \$16 \$1564 \$1121 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$30302 \$16 \$1564 \$1272 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$30304 \$153 \$1586 \$1340 \$63 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30305 \$16 \$1564 \$1303 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$30306 \$16 \$1564 \$1600 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$30308 \$16 \$1543 \$16 \$153 \$1341 VNB sky130_fd_sc_hd__inv_1
X$30309 \$153 \$1586 \$57 \$1341 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30311 \$153 \$1618 \$1340 \$509 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30313 \$153 \$1588 \$1565 \$309 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30315 \$153 \$1619 \$398 \$1651 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30316 \$153 \$1588 \$703 \$1651 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30318 \$153 \$1589 \$23 \$1651 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30319 \$153 \$1490 \$1565 \$63 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30320 \$153 \$1620 \$393 \$1651 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30322 \$16 \$149 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30324 \$16 \$509 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30325 \$16 \$1062 \$16 \$153 \$1601 VNB sky130_fd_sc_hd__clkbuf_2
X$30326 \$153 \$1619 \$1565 \$149 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30327 \$153 \$1621 \$57 \$1491 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30328 \$153 \$1621 \$1622 \$63 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30329 \$16 \$310 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30330 \$16 \$63 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30331 \$16 \$309 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30332 \$16 \$265 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30334 \$16 \$901 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30335 \$16 \$1566 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30336 \$16 \$1601 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30337 \$16 \$1566 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30338 \$16 \$1628 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30339 \$16 \$149 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30340 \$153 \$1477 \$1622 \$149 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30341 \$153 \$1534 \$23 \$1491 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30342 \$16 \$1708 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30345 \$153 \$1652 \$393 \$1491 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30346 \$16 \$1647 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30347 \$16 \$1518 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30348 \$16 \$509 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30350 \$153 \$1590 \$1342 \$509 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30351 \$16 \$309 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30352 \$153 \$1654 \$1342 \$309 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30355 \$153 \$1653 \$393 \$1255 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30356 \$153 \$1519 \$57 \$1255 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30358 \$153 \$1654 \$703 \$1255 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30359 \$16 \$309 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30360 \$16 \$178 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30361 \$153 \$1591 \$1302 \$178 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30362 \$153 \$1590 \$371 \$1255 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30366 \$153 \$1592 \$1302 \$309 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30367 \$153 \$1591 \$549 \$1343 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30369 \$16 \$63 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30370 \$153 \$1567 \$1492 \$63 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30372 \$153 \$1567 \$57 \$1414 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30374 \$16 \$1601 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30375 \$16 \$1649 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30376 \$16 \$1593 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30377 \$16 \$1599 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30378 \$16 \$149 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30379 \$153 \$1493 \$1492 \$149 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30380 \$153 \$1602 \$23 \$1414 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30381 \$16 \$1475 \$1601 \$1655 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$30383 \$16 \$1601 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30385 \$16 \$309 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30386 \$153 \$1386 \$1568 \$63 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30387 \$153 \$1387 \$1568 \$309 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30388 \$16 \$1475 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30389 \$153 \$1623 \$371 \$1414 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30390 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$30391 \$16 \$149 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30393 \$153 \$1569 \$1568 \$149 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30394 \$153 \$1668 \$371 \$1415 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30396 \$153 \$1545 \$1568 \$310 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30398 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$30399 \$153 \$1624 \$23 \$1344 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30400 \$153 \$1545 \$223 \$1344 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30401 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$30402 \$153 \$1569 \$398 \$1344 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30403 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$30404 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$30407 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$30409 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$30410 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$30411 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$30412 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$30415 \$153 \$10328 \$10554 \$10427 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30416 \$153 \$10206 \$10554 \$10368 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30417 \$16 \$10368 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30418 \$153 \$10531 \$10327 \$10511 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30419 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$30421 \$16 \$10427 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30422 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$30423 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$30425 \$153 \$10086 \$10554 \$10646 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30426 \$153 \$10207 \$10554 \$10367 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30427 \$16 \$10646 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30428 \$16 \$10367 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30429 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$30430 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$30433 \$153 \$10183 \$10554 \$10476 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30434 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$30436 \$153 \$10411 \$10705 \$10245 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30437 \$16 \$10730 \$16 \$153 \$10006 VNB sky130_fd_sc_hd__inv_1
X$30438 \$16 \$10476 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30439 \$16 \$10226 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30440 \$153 \$10593 \$10276 \$10599 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30441 \$16 \$10603 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30443 \$153 \$10302 \$10250 \$10367 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30445 \$16 \$10730 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30446 \$16 \$10730 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30447 \$153 \$10618 \$10594 \$10200 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30448 \$153 \$10428 \$10327 \$10210 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30449 \$16 \$10367 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30450 \$16 \$10200 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30451 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$30453 \$153 \$10569 \$10594 \$10368 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30454 \$16 \$10539 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30457 \$16 \$10539 \$10468 \$10512 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$30458 \$153 \$10250 \$10522 \$10512 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$30459 \$153 \$10569 \$10303 \$10599 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30460 \$16 \$10522 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30461 \$16 \$10368 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30463 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$30464 \$153 \$10533 \$10532 \$10226 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30466 \$153 \$10619 \$10532 \$10368 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30467 \$153 \$10251 \$10523 \$10469 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$30469 \$153 \$10570 \$10532 \$10646 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30470 \$16 \$10226 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30472 \$16 \$10453 \$16 \$153 \$10211 VNB sky130_fd_sc_hd__inv_1
X$30474 \$153 \$10534 \$10259 \$10476 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30475 \$153 \$10429 \$10705 \$10211 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30476 \$153 \$10570 \$10318 \$10745 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30477 \$16 \$10476 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30478 \$16 \$10453 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30479 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$30480 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$30481 \$16 \$10555 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30482 \$153 \$10489 \$10259 \$10367 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30484 \$153 \$10534 \$10705 \$10246 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30486 \$16 \$10555 \$16 \$153 \$10246 VNB sky130_fd_sc_hd__inv_1
X$30487 \$153 \$9897 \$8737 \$9866 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30488 \$153 \$10489 \$10330 \$10246 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30489 \$153 \$10620 \$10199 \$10476 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30490 \$16 \$10427 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30491 \$16 \$10367 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30493 \$153 \$10535 \$10199 \$10367 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30494 \$153 \$10535 \$10330 \$10212 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30495 \$153 \$10490 \$10318 \$10212 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30496 \$153 \$10092 \$8726 \$9866 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30497 \$153 \$10491 \$10524 \$10295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30499 \$153 \$10571 \$10524 \$10368 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30500 \$153 \$10491 \$10276 \$10513 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30501 \$153 \$10571 \$10303 \$10513 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30502 \$16 \$10368 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30504 \$16 \$10367 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30507 \$153 \$10536 \$10252 \$10367 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30509 \$16 \$10427 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30510 \$16 \$10476 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30512 \$153 \$10431 \$10705 \$10331 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30513 \$153 \$10600 \$10318 \$10513 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30514 \$153 \$10536 \$10330 \$10331 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30515 \$16 \$10621 \$16 \$153 \$10331 VNB sky130_fd_sc_hd__inv_1
X$30517 \$16 \$10367 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30518 \$153 \$10492 \$10456 \$10367 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30519 \$16 \$10621 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30521 \$16 \$10621 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30523 \$16 \$6647 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30524 \$153 \$10432 \$10161 \$10334 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30526 \$153 \$10492 \$10330 \$10334 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30527 \$153 \$6647 \$9339 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$30528 \$16 \$10226 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30531 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$30532 \$153 \$10493 \$10456 \$10200 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30533 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$30534 \$153 \$10601 \$10318 \$10334 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30535 \$153 \$10493 \$10088 \$10334 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30536 \$16 \$10705 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30537 \$16 \$10295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30540 \$153 \$153 \$10705 \$10602 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30541 \$16 \$10200 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30542 \$16 \$6712 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30543 \$153 \$6712 \$9869 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$30545 \$153 \$153 \$10276 \$10602 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30546 \$153 \$10320 \$10603 \$10537 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$30549 \$16 \$10348 \$10525 \$10537 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$30550 \$16 \$10348 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30551 \$16 \$10603 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30552 \$153 \$10556 \$10320 \$10514 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30553 \$153 \$10457 \$10320 \$10526 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30554 \$153 \$10458 \$10320 \$10605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30555 \$16 \$10526 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30556 \$16 \$10514 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30559 \$16 \$10202 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30560 \$16 \$10145 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30561 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$30562 \$153 \$10557 \$10653 \$10338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30563 \$153 \$10556 \$10538 \$10369 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30564 \$16 \$10605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30565 \$16 \$10147 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30566 \$16 \$10338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30567 \$153 \$10622 \$10653 \$10298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30570 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$30571 \$16 \$10539 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30572 \$153 \$10494 \$10247 \$10369 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30573 \$153 \$10557 \$10309 \$10477 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30574 \$16 \$10298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30576 \$153 \$10336 \$10400 \$10382 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30577 \$16 \$10539 \$10525 \$10623 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$30578 \$16 \$10522 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30581 \$153 \$10572 \$10400 \$10526 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30583 \$153 \$10540 \$10400 \$10605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30584 \$153 \$10572 \$10516 \$10337 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30585 \$16 \$10526 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30586 \$16 \$10382 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30587 \$153 \$10604 \$10538 \$10337 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30590 \$153 \$10380 \$10523 \$10541 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$30591 \$153 \$10307 \$10247 \$10337 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30592 \$153 \$10542 \$10380 \$10514 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30593 \$16 \$10523 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30595 \$153 \$10496 \$10247 \$10339 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30597 \$153 \$10495 \$10344 \$10339 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30598 \$153 \$10542 \$10538 \$10339 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30599 \$16 \$10514 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30601 \$153 \$10573 \$10380 \$10605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30602 \$153 \$10497 \$10380 \$10526 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30604 \$153 \$10573 \$10686 \$10339 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30605 \$153 \$10497 \$10516 \$10339 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30607 \$153 \$10543 \$10381 \$10526 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30608 \$16 \$10526 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30610 \$153 \$10498 \$10344 \$10515 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30611 \$153 \$10543 \$10516 \$10515 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30612 \$16 \$10555 \$16 \$153 \$10515 VNB sky130_fd_sc_hd__inv_1
X$30614 \$16 \$10526 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30615 \$153 \$10499 \$10381 \$10470 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30616 \$16 \$10605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30617 \$153 \$10544 \$10381 \$10514 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30618 \$153 \$10544 \$10538 \$10515 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30619 \$16 \$10514 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30620 \$16 \$10621 \$16 \$153 \$10249 VNB sky130_fd_sc_hd__inv_1
X$30621 \$153 \$10574 \$10340 \$10526 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30624 \$153 \$10435 \$10098 \$10515 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30625 \$153 \$10499 \$10247 \$10515 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30626 \$153 \$10574 \$10516 \$10249 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30627 \$153 \$10545 \$10344 \$10249 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30628 \$16 \$10526 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30629 \$16 \$10606 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30630 \$16 \$10624 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30631 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$30633 \$153 \$10625 \$10340 \$10605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30634 \$153 \$10546 \$10538 \$10249 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30635 \$153 \$10403 \$10323 \$10470 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30637 \$153 \$10547 \$10323 \$10526 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30639 \$16 \$10470 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30641 \$153 \$10547 \$10516 \$10343 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30642 \$16 \$10526 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30643 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$30644 \$153 \$10575 \$10607 \$10514 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30645 \$16 \$10514 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30647 \$16 \$9845 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30648 \$153 \$10205 \$10606 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$30651 \$153 \$10575 \$10538 \$10608 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30652 \$16 \$10205 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30653 \$153 \$10558 \$10607 \$10470 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30654 \$153 \$10576 \$10607 \$10338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30657 \$153 \$10576 \$10309 \$10608 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30658 \$16 \$10139 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30659 \$16 \$7934 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30660 \$153 \$10527 \$10605 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$30661 \$153 \$10408 \$10526 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$30662 \$153 \$10265 \$8340 \$10538 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30664 \$153 \$9339 \$10735 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$30665 \$16 \$7934 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30666 \$153 \$9228 \$9133 \$7994 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30668 \$153 \$10610 \$10714 \$10609 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30669 \$16 \$10238 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30670 \$16 \$10527 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30673 \$16 \$9227 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30674 \$16 \$9869 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30675 \$153 \$9869 \$10611 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$30677 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30678 \$153 \$10145 \$8340 \$10714 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30679 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30680 \$153 \$10319 \$8340 \$10417 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30681 \$16 \$10686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30682 \$16 \$9275 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30684 \$153 \$6921 \$8320 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$30685 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30687 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30688 \$16 \$16 \$153 VNB sky130_fd_sc_hd__conb_1
X$30689 \$153 \$153 \$10472 \$10479 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30690 \$16 \$6921 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30692 \$16 \$10478 \$16 \$153 \$10479 VNB sky130_fd_sc_hd__clkbuf_2
X$30693 \$153 \$153 \$10471 \$10479 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30695 \$153 \$153 \$10370 \$10479 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30696 \$16 \$10370 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30697 \$153 \$153 \$10417 \$10479 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30698 \$16 \$10300 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30699 \$153 \$10549 \$10463 \$10300 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30700 \$153 \$10464 \$10463 \$10578 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30702 \$153 \$10612 \$10501 \$10480 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30703 \$16 \$10714 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30704 \$16 \$10478 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30705 \$153 \$10613 \$10471 \$10372 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30706 \$16 \$10473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30707 \$153 \$10465 \$10463 \$10473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30708 \$153 \$10713 \$10919 \$10372 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30709 \$153 \$10596 \$10714 \$10372 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30711 \$153 \$10549 \$10417 \$10372 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30712 \$153 \$10577 \$10528 \$10551 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30713 \$153 \$10481 \$10528 \$10300 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30714 \$16 \$10551 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30715 \$153 \$10550 \$10528 \$10473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30718 \$153 \$10577 \$10471 \$10482 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30719 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$30720 \$153 \$10437 \$10472 \$10482 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30722 \$16 \$10578 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30723 \$153 \$10579 \$10474 \$10578 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30724 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$30725 \$16 \$10386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30727 \$153 \$10483 \$10474 \$10386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30728 \$153 \$10614 \$10833 \$10372 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30729 \$153 \$10579 \$10370 \$10373 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30730 \$153 \$10502 \$10474 \$10473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30731 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$30732 \$16 \$10300 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30734 \$153 \$10559 \$10404 \$10300 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30735 \$153 \$10503 \$10404 \$10473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30737 \$153 \$10580 \$10404 \$10551 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30738 \$16 \$10551 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30740 \$16 \$10552 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30741 \$16 \$10611 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30743 \$153 \$9974 \$8917 \$9642 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30745 \$16 \$10551 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30746 \$153 \$10581 \$10387 \$10551 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30747 \$16 \$9642 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30749 \$153 \$10553 \$10387 \$10611 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30750 \$16 \$10615 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30751 \$16 \$10597 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30752 \$153 \$9975 \$8676 \$9642 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30754 \$16 \$10735 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30755 \$153 \$10582 \$10387 \$10735 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30756 \$153 \$10406 \$10370 \$10374 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30757 \$153 \$10407 \$10472 \$10374 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30758 \$16 \$10597 \$16 \$153 \$10374 VNB sky130_fd_sc_hd__inv_1
X$30760 \$153 \$10583 \$10475 \$10735 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30763 \$153 \$10504 \$10475 \$10386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30764 \$153 \$10440 \$10501 \$10374 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30765 \$153 \$10441 \$10417 \$10517 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30766 \$153 \$10583 \$10919 \$10517 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30767 \$16 \$10578 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30768 \$153 \$10505 \$10388 \$10578 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30770 \$153 \$10584 \$10388 \$10611 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30771 \$153 \$10505 \$10370 \$10375 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30773 \$16 \$10735 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30774 \$153 \$10585 \$10388 \$10735 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30775 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$30777 \$153 \$10443 \$10472 \$10375 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30779 \$16 \$10551 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30781 \$153 \$10586 \$10388 \$10551 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30782 \$16 \$10809 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30784 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30785 \$153 \$10390 \$8340 \$10815 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30786 \$16 \$10815 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30788 \$153 \$10586 \$10471 \$10375 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30789 \$16 \$10529 \$16 \$153 \$10375 VNB sky130_fd_sc_hd__inv_1
X$30790 \$153 \$10316 \$8340 \$10642 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30791 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30792 \$153 \$10158 \$8340 \$10466 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30793 \$16 \$16 \$153 VNB sky130_fd_sc_hd__conb_1
X$30795 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30796 \$153 \$10268 \$8340 \$10587 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30798 \$16 \$10642 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30799 \$16 \$10560 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30800 \$16 \$10376 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30801 \$16 \$10466 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30803 \$16 \$10694 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30804 \$153 \$10408 \$10564 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$30805 \$16 \$10587 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30806 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$30807 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$30810 \$16 \$11068 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30811 \$153 \$6994 \$10408 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$30812 \$153 \$10485 \$10616 \$10326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30814 \$153 \$10588 \$10587 \$10484 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30815 \$16 \$6994 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30816 \$16 \$10326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30819 \$153 \$10561 \$10616 \$10346 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30820 \$153 \$10598 \$10616 \$10446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30821 \$16 \$10139 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30822 \$153 \$10561 \$10285 \$10484 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30823 \$153 \$10139 \$10617 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$30824 \$16 \$10346 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30826 \$153 \$10598 \$10376 \$10484 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30827 \$153 \$10486 \$10285 \$11016 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30828 \$153 \$10562 \$10530 \$10393 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30829 \$153 \$10562 \$10694 \$10518 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30830 \$16 \$10393 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30831 \$16 \$10446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30833 \$16 \$10392 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30835 \$16 \$10467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30836 \$153 \$10506 \$10530 \$10346 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30837 \$153 \$10589 \$10530 \$10467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30839 \$153 \$10563 \$10444 \$10326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30840 \$16 \$10346 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30841 \$16 \$10326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30842 \$16 \$10897 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30843 \$16 \$10392 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30846 \$16 \$10617 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30847 \$153 \$10626 \$10444 \$10617 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30848 \$153 \$10506 \$10285 \$10518 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30850 \$153 \$10507 \$10694 \$10519 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30851 \$153 \$10589 \$10587 \$10518 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30852 \$16 \$10446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30854 \$153 \$10563 \$10466 \$10519 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30855 \$153 \$10487 \$10444 \$10446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30857 \$16 \$10467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30858 \$153 \$10627 \$10394 \$10467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30859 \$16 \$10346 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30860 \$16 \$10393 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30861 \$153 \$10508 \$10394 \$10393 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30863 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$30864 \$16 \$10564 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30865 \$153 \$10590 \$10394 \$10564 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30866 \$16 \$10446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30867 \$153 \$10508 \$10694 \$10520 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30868 \$153 \$10509 \$10376 \$10520 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30869 \$153 \$10590 \$10642 \$10520 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30872 \$16 \$10392 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30873 \$153 \$10565 \$10395 \$10392 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30874 \$16 \$10564 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30875 \$153 \$10628 \$10395 \$10564 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30876 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$30877 \$16 \$10661 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30878 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$30880 \$153 \$10449 \$10376 \$10521 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30883 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$30884 \$16 \$10617 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30885 \$153 \$10566 \$10325 \$10393 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30886 \$153 \$10629 \$10325 \$10617 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30888 \$16 \$10597 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30889 \$16 \$10222 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30890 \$16 \$10467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30891 \$153 \$9709 \$8965 \$10222 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30893 \$16 \$8429 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30894 \$153 \$8878 \$7375 \$8429 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30895 \$153 \$10591 \$10396 \$10467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30896 \$153 \$9381 \$7180 \$8429 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30897 \$153 \$9943 \$9256 \$10510 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30898 \$16 \$10409 \$10644 \$10630 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$30900 \$16 \$8429 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30901 \$153 \$9645 \$9122 \$9646 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30902 \$153 \$10631 \$10396 \$10564 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30903 \$153 \$10365 \$8923 \$10112 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30904 \$153 \$8055 \$7607 \$7076 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30905 \$16 \$7076 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30906 \$16 \$10564 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30907 \$153 \$9710 \$8996 \$9646 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30909 \$153 \$10567 \$10397 \$10393 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30910 \$153 \$10632 \$10592 \$10564 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30911 \$153 \$10292 \$9122 \$10112 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30912 \$153 \$9712 \$8923 \$9646 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30913 \$16 \$10393 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30914 \$16 \$10446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30916 \$153 \$10633 \$10592 \$10446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30917 \$16 \$10617 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30918 \$153 \$10568 \$10397 \$10617 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30919 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$30920 \$153 \$9784 \$9103 \$9646 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30921 \$153 \$9714 \$8965 \$9646 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30923 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$30924 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$30925 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$30926 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$30927 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$30928 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$30930 \$153 \$7919 \$7864 \$6981 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30931 \$153 \$8000 \$7864 \$6783 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30932 \$153 \$7920 \$7864 \$6784 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30933 \$153 \$8000 \$6749 \$7765 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30935 \$153 \$7794 \$7864 \$6907 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30936 \$153 \$7920 \$6794 \$7765 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30937 \$153 \$7883 \$6732 \$7765 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30938 \$16 \$6907 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30940 \$16 \$7816 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30941 \$16 \$8001 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30942 \$16 \$6784 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30943 \$153 \$8033 \$6732 \$8034 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30944 \$16 \$6987 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30946 \$153 \$7795 \$7864 \$6979 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30948 \$16 \$8001 \$16 \$153 \$7765 VNB sky130_fd_sc_hd__inv_1
X$30949 \$153 \$7864 \$7884 \$8002 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$30950 \$16 \$6979 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30951 \$153 \$7796 \$7784 \$6979 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30952 \$16 \$8001 \$8024 \$8002 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$30955 \$153 \$7940 \$7784 \$7041 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30957 \$153 \$7940 \$6996 \$7711 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30958 \$153 \$7941 \$6749 \$7711 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30959 \$16 \$7041 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30960 \$16 \$8003 \$16 \$153 \$7711 VNB sky130_fd_sc_hd__inv_1
X$30961 \$153 \$7784 \$8438 \$8056 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$30962 \$16 \$6979 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30966 \$16 \$6981 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30967 \$16 \$8003 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30968 \$16 \$8438 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30969 \$153 \$7921 \$7620 \$6979 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30970 \$153 \$7865 \$7620 \$6860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30971 \$16 \$6979 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30972 \$153 \$7921 \$6995 \$7587 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30973 \$16 \$6860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30976 \$153 \$8035 \$6719 \$8036 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30977 \$153 \$7961 \$7620 \$6981 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30978 \$153 \$7620 \$7655 \$7962 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$30979 \$16 \$7922 \$8024 \$7962 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$30980 \$153 \$7885 \$6719 \$7587 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30981 \$16 \$7922 \$16 \$153 \$7587 VNB sky130_fd_sc_hd__inv_1
X$30983 \$16 \$6981 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30985 \$16 \$6860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30986 \$153 \$8057 \$7866 \$7041 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30987 \$153 \$7963 \$7866 \$6792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$30989 \$16 \$6792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30990 \$153 \$6912 \$6995 \$6733 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30991 \$16 \$7041 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30992 \$16 \$6784 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30995 \$16 \$6733 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30996 \$153 \$7621 \$6749 \$7608 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$30997 \$16 \$6733 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30998 \$16 \$6912 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$30999 \$16 \$7816 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31000 \$153 \$7987 \$7866 \$6783 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31001 \$16 \$6863 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31002 \$16 \$7135 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31003 \$153 \$7818 \$6794 \$7608 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31005 \$16 \$6783 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31006 \$153 \$7817 \$6732 \$7608 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31009 \$16 \$7040 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31011 \$153 \$7964 \$7701 \$6981 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31012 \$153 \$7988 \$7701 \$6907 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31013 \$153 \$7965 \$7701 \$6784 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31014 \$16 \$6981 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31015 \$16 \$6907 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31016 \$16 \$7887 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31019 \$153 \$8057 \$6996 \$7609 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31020 \$153 \$7932 \$6930 \$7609 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31021 \$153 \$8004 \$6794 \$7609 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31022 \$153 \$7886 \$6995 \$7609 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31024 \$153 \$8058 \$7703 \$7041 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31026 \$16 \$6979 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31029 \$16 \$6981 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31031 \$153 \$7966 \$6719 \$7768 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31032 \$16 \$7041 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31034 \$16 \$6783 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31035 \$153 \$8059 \$7703 \$6783 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31036 \$153 \$7942 \$6732 \$7768 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31038 \$16 \$6753 \$8195 \$7943 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$31039 \$153 \$7337 \$6903 \$7943 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$31041 \$16 \$8125 \$8195 \$8060 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$31042 \$16 \$8125 \$16 \$153 \$7768 VNB sky130_fd_sc_hd__inv_1
X$31043 \$153 \$8062 \$7989 \$8037 \$8026 \$8005 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$31044 \$16 \$6981 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31046 \$153 \$7714 \$7705 \$7770 \$7771 \$7785 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$31047 \$153 \$8063 \$7989 \$8026 \$8005 \$8037 \$16 \$16 VNB
+ sky130_fd_sc_hd__nor4b_2
X$31050 \$153 \$7848 \$6749 \$7772 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31051 \$153 \$8064 \$8005 \$8037 \$8026 \$7989 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$31052 \$153 \$7964 \$6930 \$7772 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31053 \$153 \$8026 \$7989 \$8065 \$8005 \$8037 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$31054 \$16 \$7770 \$7705 \$7771 \$7785 \$16 \$153 \$7713 VNB
+ sky130_fd_sc_hd__and4_2
X$31055 \$16 \$7944 \$16 \$153 \$7705 VNB sky130_fd_sc_hd__clkbuf_2
X$31056 \$16 \$7945 \$8061 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$31057 \$16 \$7889 \$16 \$153 \$7771 VNB sky130_fd_sc_hd__clkbuf_2
X$31059 \$16 \$7967 \$16 \$153 \$7770 VNB sky130_fd_sc_hd__clkbuf_2
X$31060 \$16 \$7944 \$16 \$153 \$7470 VNB sky130_fd_sc_hd__clkbuf_2
X$31061 \$16 \$7786 \$16 \$153 \$8038 VNB sky130_fd_sc_hd__clkbuf_2
X$31063 \$16 \$7559 \$16 \$153 \$7889 VNB sky130_fd_sc_hd__clkbuf_2
X$31064 \$16 \$7889 \$16 \$153 \$8066 VNB sky130_fd_sc_hd__clkbuf_2
X$31065 \$16 \$6540 \$16 \$153 \$7944 VNB sky130_fd_sc_hd__clkbuf_2
X$31066 \$16 \$7944 \$16 \$153 \$8067 VNB sky130_fd_sc_hd__clkbuf_2
X$31067 \$16 \$7945 \$8119 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$31069 \$16 \$8039 \$16 \$153 \$8003 VNB sky130_fd_sc_hd__clkbuf_2
X$31070 \$16 \$7867 \$7800 \$7859 \$153 \$7967 \$16 VNB sky130_fd_sc_hd__and3b_4
X$31071 \$16 \$7559 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31072 \$153 \$7624 \$7655 \$8068 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$31074 \$16 \$7867 \$7859 \$7800 \$153 \$16 \$7891 VNB sky130_fd_sc_hd__and3_4
X$31075 \$16 \$7890 \$16 \$153 \$7990 VNB sky130_fd_sc_hd__clkbuf_2
X$31076 \$16 \$6540 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31078 \$153 \$7868 \$7946 \$6862 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31079 \$16 \$7922 \$16 \$153 \$7611 VNB sky130_fd_sc_hd__inv_1
X$31080 \$153 \$7969 \$7946 \$6754 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31083 \$153 \$7969 \$6756 \$7787 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31084 \$16 \$5477 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31085 \$16 \$6451 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31087 \$153 \$7970 \$7946 \$6916 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31088 \$153 \$8069 \$7946 \$7060 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31089 \$16 \$6754 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31090 \$153 \$7970 \$6867 \$7787 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31093 \$153 \$7869 \$7624 \$7060 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31094 \$16 \$6916 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31095 \$16 \$8003 \$7968 \$8006 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$31096 \$153 \$7627 \$8438 \$8006 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$31097 \$16 \$7060 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31098 \$16 \$8001 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31099 \$16 \$8438 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31100 \$16 \$6916 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31101 \$153 \$7892 \$7627 \$6916 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31103 \$16 \$8003 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31104 \$153 \$8007 \$7627 \$6862 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31105 \$153 \$7870 \$7627 \$6771 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31106 \$153 \$8007 \$7003 \$7562 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31108 \$16 \$6862 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31109 \$16 \$6771 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31112 \$153 \$7991 \$7947 \$7044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31113 \$153 \$7971 \$7947 \$6991 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31114 \$153 \$7971 \$6992 \$8040 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31115 \$16 \$7548 \$16 \$153 \$7968 VNB sky130_fd_sc_hd__clkbuf_2
X$31116 \$153 \$7972 \$7947 \$6797 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31119 \$16 \$6991 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31120 \$16 \$6916 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31121 \$16 \$7044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31122 \$153 \$7972 \$6906 \$8040 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31123 \$153 \$7991 \$7006 \$8040 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31124 \$153 \$8070 \$7707 \$7044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31125 \$16 \$6797 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31127 \$16 \$7973 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31128 \$16 \$8177 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31130 \$16 \$7548 \$16 \$153 \$7804 VNB sky130_fd_sc_hd__clkbuf_2
X$31131 \$153 \$7893 \$6324 \$7718 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31132 \$153 \$7746 \$6906 \$7718 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31133 \$16 \$7044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31134 \$16 \$6754 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31135 \$16 \$7973 \$7804 \$8008 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$31136 \$153 \$7974 \$7684 \$6771 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31137 \$153 \$7825 \$7006 \$7895 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31139 \$153 \$8041 \$6992 \$7895 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31140 \$153 \$7974 \$6865 \$7895 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31141 \$153 \$8071 \$7684 \$6916 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31142 \$16 \$6771 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31143 \$16 \$7992 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31144 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$31145 \$153 \$7896 \$6906 \$7895 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31146 \$16 \$6916 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31149 \$153 \$7826 \$6756 \$7895 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31150 \$16 \$7992 \$16 \$153 \$7720 VNB sky130_fd_sc_hd__inv_1
X$31151 \$153 \$8009 \$7788 \$6991 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31152 \$153 \$7975 \$6324 \$7895 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31153 \$153 \$7747 \$7003 \$7895 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31154 \$153 \$8009 \$6992 \$7720 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31155 \$153 \$7774 \$6906 \$7720 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31157 \$153 \$8010 \$7788 \$6771 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31158 \$153 \$7479 \$7887 \$7948 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$31159 \$153 \$8010 \$6865 \$7720 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31160 \$16 \$7663 \$7804 \$7948 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$31161 \$16 \$6753 \$7804 \$7899 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$31164 \$153 \$7897 \$6865 \$7612 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31165 \$153 \$8011 \$8027 \$6991 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31166 \$153 \$7708 \$6887 \$7828 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$31167 \$153 \$8011 \$6992 \$7933 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31168 \$16 \$6991 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31170 \$153 \$7923 \$8027 \$7060 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31173 \$16 \$6887 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31175 \$153 \$8042 \$7003 \$7933 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31176 \$153 \$8012 \$8027 \$6771 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31177 \$153 \$7923 \$6324 \$7933 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31178 \$16 \$6916 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31179 \$16 \$7060 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31182 \$16 \$7934 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31183 \$153 \$8012 \$6865 \$7933 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31184 \$16 \$7949 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31185 \$16 \$7949 \$7829 \$7934 \$153 \$7288 \$16 VNB sky130_fd_sc_hd__and3b_4
X$31186 \$16 \$6771 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31188 \$153 \$153 \$6756 \$7872 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31189 \$153 \$153 \$6324 \$7872 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31190 \$16 \$16 \$153 VNB sky130_fd_sc_hd__conb_1
X$31191 \$16 \$7288 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31192 \$16 \$6771 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31194 \$16 \$7829 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31197 \$153 \$153 \$6865 \$7872 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31198 \$153 \$153 \$6906 \$7872 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31200 \$153 \$153 \$7006 \$7872 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31201 \$153 \$7775 \$7215 \$7296 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31202 \$153 \$7900 \$7490 \$7296 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31203 \$153 \$8072 \$8028 \$7387 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31205 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$31206 \$16 \$7082 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31208 \$153 \$7873 \$8028 \$7082 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31209 \$153 \$7993 \$8028 \$7328 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31210 \$16 \$7793 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31211 \$16 \$7328 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31212 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$31214 \$16 \$7793 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31215 \$16 \$7445 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31217 \$16 \$7029 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31218 \$153 \$7977 \$7874 \$7445 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31219 \$153 \$7935 \$7874 \$7029 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31221 \$153 \$7935 \$7066 \$7924 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31222 \$153 \$7977 \$7327 \$7924 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31223 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$31225 \$153 \$7902 \$7215 \$7924 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31226 \$16 \$7328 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31227 \$153 \$7950 \$7874 \$7328 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31228 \$153 \$7666 \$7065 \$7597 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31229 \$153 \$7950 \$7366 \$7924 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31231 \$16 \$9150 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31232 \$16 \$7129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31233 \$16 \$7067 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31234 \$16 \$7445 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31236 \$153 \$7925 \$7876 \$7445 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31237 \$153 \$8013 \$7876 \$7129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31238 \$16 \$7994 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31239 \$153 \$7925 \$7327 \$7789 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31241 \$16 \$8073 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31242 \$16 \$7387 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31243 \$153 \$8074 \$7876 \$7387 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31244 \$16 \$7082 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31246 \$16 \$7995 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31247 \$16 \$7239 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31248 \$153 \$7978 \$7876 \$7239 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31249 \$153 \$8014 \$7215 \$8043 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31250 \$16 \$7029 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31251 \$153 \$7979 \$7635 \$7029 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31252 \$16 \$7994 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31253 \$16 \$8044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31254 \$16 \$7996 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31256 \$153 \$7978 \$7482 \$7789 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31257 \$153 \$7878 \$7635 \$7067 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31259 \$153 \$7979 \$7066 \$7571 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31260 \$153 \$8045 \$7366 \$7571 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31261 \$16 \$7067 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31262 \$16 \$7129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31264 \$153 \$7997 \$8029 \$7129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31265 \$153 \$7905 \$7327 \$7571 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31266 \$153 \$7980 \$7636 \$7129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31267 \$16 \$7129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31269 \$153 \$8046 \$7066 \$8222 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31270 \$153 \$7906 \$7366 \$7613 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31272 \$153 \$7980 \$7215 \$7613 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31273 \$16 \$7691 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31274 \$16 \$7952 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31275 \$16 \$7691 \$16 \$153 \$7613 VNB sky130_fd_sc_hd__inv_1
X$31277 \$153 \$8015 \$7065 \$8047 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31278 \$153 \$7907 \$7482 \$7613 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31279 \$153 \$7636 \$7915 \$7836 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$31281 \$16 \$7952 \$7673 \$7951 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$31284 \$153 \$7790 \$8772 \$7951 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$31286 \$16 \$7445 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31287 \$153 \$8075 \$7790 \$7445 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31288 \$16 \$8772 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31289 \$16 \$7328 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31290 \$153 \$7981 \$7790 \$7328 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31291 \$16 \$7129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31292 \$16 \$7082 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31294 \$153 \$8076 \$8030 \$7082 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31295 \$153 \$7998 \$7790 \$7129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31296 \$153 \$7981 \$7366 \$7726 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31297 \$16 \$7952 \$16 \$153 \$7726 VNB sky130_fd_sc_hd__inv_1
X$31299 \$16 \$7328 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31300 \$16 \$7029 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31304 \$153 \$8016 \$7953 \$7082 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31305 \$153 \$7982 \$7953 \$7328 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31306 \$16 \$7952 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31307 \$153 \$7982 \$7366 \$8048 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31308 \$153 \$7687 \$7215 \$7728 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31309 \$16 \$7067 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31311 \$153 \$7926 \$7953 \$7067 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31312 \$153 \$8016 \$7065 \$8048 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31314 \$16 \$7445 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31315 \$153 \$7983 \$7953 \$7445 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31316 \$153 \$7926 \$6582 \$8048 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31318 \$16 \$7793 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31320 \$153 \$7983 \$7327 \$8048 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31321 \$16 \$7239 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31323 \$16 \$8049 \$16 \$153 \$7881 VNB sky130_fd_sc_hd__clkbuf_2
X$31324 \$16 \$8051 \$16 \$153 \$7791 VNB sky130_fd_sc_hd__clkbuf_2
X$31325 \$16 \$7793 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31326 \$153 \$8077 \$7881 \$7880 \$7791 \$7792 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$31327 \$153 \$7729 \$7792 \$7880 \$7881 \$7791 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$31328 \$16 \$6540 \$16 \$153 \$8050 VNB sky130_fd_sc_hd__clkbuf_2
X$31329 \$153 \$7881 \$7791 \$7730 \$7792 \$7880 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$31330 \$16 \$6540 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31333 \$16 \$8078 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31334 \$153 \$7881 \$7792 \$7641 \$7791 \$7880 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$31335 \$16 \$7984 \$16 \$153 \$7130 VNB sky130_fd_sc_hd__clkbuf_2
X$31336 \$16 \$7927 \$7954 \$7936 \$7955 \$16 \$153 \$7999 VNB
+ sky130_fd_sc_hd__and4_2
X$31338 \$16 \$7377 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31339 \$153 \$7984 \$7955 \$7927 \$7936 \$7954 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$31340 \$153 \$7908 \$7936 \$7927 \$7955 \$7954 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$31341 \$16 \$8049 \$16 \$153 \$7936 VNB sky130_fd_sc_hd__clkbuf_2
X$31342 \$16 \$8051 \$16 \$153 \$7955 VNB sky130_fd_sc_hd__clkbuf_2
X$31344 \$153 \$8017 \$7955 \$7936 \$7954 \$7927 \$16 \$16 VNB
+ sky130_fd_sc_hd__nor4b_2
X$31345 \$153 \$7780 \$7954 \$7927 \$7936 \$7955 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$31346 \$153 \$7936 \$7954 \$7909 \$7955 \$7927 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$31347 \$153 \$7936 \$7955 \$8052 \$7954 \$7927 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$31348 \$16 \$7133 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31349 \$16 \$8017 \$16 \$153 \$7495 VNB sky130_fd_sc_hd__clkbuf_2
X$31350 \$153 \$7910 \$7462 \$7731 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31351 \$16 \$16 \$153 VNB sky130_fd_sc_hd__conb_1
X$31353 \$153 \$153 \$7462 \$8186 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31354 \$153 \$7937 \$7642 \$7133 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31356 \$153 \$7911 \$7375 \$7731 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31358 \$153 \$7937 \$7180 \$7731 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31359 \$153 \$8080 \$8018 \$7464 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31361 \$16 \$7133 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31362 \$16 \$7307 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31363 \$153 \$7938 \$7208 \$7928 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31364 \$16 \$7464 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31366 \$16 \$7353 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31367 \$153 \$8019 \$8018 \$7307 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31368 \$153 \$7929 \$8018 \$7377 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31370 \$153 \$7929 \$7462 \$7928 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31371 \$153 \$8019 \$7607 \$7928 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31373 \$153 \$7508 \$7208 \$7734 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31374 \$16 \$7464 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31375 \$153 \$8020 \$7862 \$7464 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31376 \$153 \$7912 \$7375 \$7734 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31378 \$153 \$7957 \$7607 \$7939 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31379 \$153 \$8020 \$7639 \$7939 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31381 \$16 \$7353 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31382 \$16 \$7174 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31383 \$153 \$8021 \$7862 \$7353 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31384 \$153 \$7930 \$7862 \$7174 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31388 \$153 \$8021 \$7375 \$7939 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31389 \$153 \$7930 \$7376 \$7939 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31390 \$153 \$7913 \$7208 \$7939 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31391 \$153 \$8053 \$7180 \$8291 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31392 \$153 \$7308 \$7208 \$6985 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31393 \$153 \$8082 \$8189 \$7131 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31395 \$16 \$7904 \$16 \$153 \$7616 VNB sky130_fd_sc_hd__inv_1
X$31396 \$16 \$7377 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31398 \$16 \$7464 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31399 \$16 \$7353 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31400 \$153 \$7931 \$7710 \$7464 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31401 \$153 \$8022 \$7710 \$7353 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31402 \$16 \$7147 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31403 \$153 \$7931 \$7639 \$7616 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31404 \$16 \$7131 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31406 \$153 \$8022 \$7375 \$7616 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31408 \$153 \$7688 \$8772 \$7958 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$31409 \$153 \$8054 \$7180 \$8098 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31410 \$153 \$7813 \$7688 \$7377 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31411 \$16 \$7952 \$7496 \$7958 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$31412 \$16 \$7952 \$16 \$153 \$7580 VNB sky130_fd_sc_hd__inv_1
X$31414 \$153 \$7914 \$7375 \$7580 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31415 \$153 \$8023 \$8031 \$7131 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31417 \$153 \$7698 \$7915 \$7959 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$31418 \$16 \$7691 \$7496 \$7959 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$31419 \$153 \$7985 \$7698 \$7353 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31422 \$153 \$8083 \$7698 \$7131 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31424 \$153 \$7841 \$7180 \$7882 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31425 \$153 \$8084 \$7698 \$7307 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31426 \$16 \$7307 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31427 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$31429 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$31431 \$16 \$8359 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31432 \$16 \$7147 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31433 \$153 \$7454 \$7639 \$7217 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31434 \$16 \$8032 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31435 \$16 \$7377 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31436 \$153 \$8085 \$7863 \$7377 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31437 \$153 \$7272 \$7863 \$7147 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31440 \$16 \$7174 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31442 \$153 \$7956 \$7863 \$7174 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31443 \$16 \$7307 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31444 \$153 \$8055 \$7863 \$7307 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31445 \$16 \$7695 \$7496 \$7814 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$31446 \$16 \$7695 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31447 \$16 \$8265 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31448 \$16 \$7353 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31451 \$16 \$7431 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31452 \$16 \$7353 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31453 \$16 \$7377 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31454 \$153 \$7069 \$7960 \$7353 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31455 \$153 \$7986 \$7647 \$7377 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31456 \$153 \$7762 \$7463 \$7782 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31457 \$16 \$7131 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31458 \$153 \$7048 \$7960 \$7131 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31460 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$31462 \$16 \$7377 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31463 \$153 \$8086 \$7960 \$7377 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31464 \$153 \$10728 \$7960 \$7174 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31465 \$153 \$7918 \$7607 \$7782 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31466 \$16 \$7174 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31468 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$31470 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$31471 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$31472 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$31473 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$31474 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$31476 \$16 \$6813 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31477 \$153 \$8855 \$8895 \$9129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31478 \$153 \$8948 \$8895 \$8580 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31480 \$153 \$8855 \$8737 \$8882 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31481 \$16 \$8580 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31483 \$153 \$8978 \$8912 \$8882 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31484 \$153 \$8799 \$8667 \$8828 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31485 \$153 \$8948 \$8194 \$8882 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31486 \$16 \$8828 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31487 \$153 \$8896 \$8885 \$8679 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31489 \$153 \$8949 \$8895 \$9026 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31491 \$16 \$9026 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31492 \$16 \$9026 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31494 \$16 \$6988 \$16 \$153 \$8882 VNB sky130_fd_sc_hd__inv_1
X$31495 \$153 \$8895 \$6888 \$8856 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$31496 \$153 \$8949 \$8726 \$8882 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31497 \$153 \$8979 \$8457 \$8679 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31498 \$153 \$8434 \$8722 \$8715 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31501 \$153 \$8435 \$8722 \$8950 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31502 \$153 \$8910 \$8722 \$8828 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31503 \$153 \$8980 \$8885 \$8883 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31504 \$16 \$8950 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31505 \$16 \$8828 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31507 \$16 \$8724 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31508 \$153 \$8909 \$8209 \$8883 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31509 \$16 \$6888 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31510 \$16 \$6988 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31511 \$153 \$8884 \$8533 \$8828 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31512 \$153 \$8827 \$8533 \$9129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31513 \$16 \$8828 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31514 \$16 \$7378 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31515 \$16 \$9129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31516 \$153 \$8780 \$8638 \$8723 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31519 \$153 \$8969 \$8457 \$8883 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31520 \$153 \$8884 \$8885 \$8723 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31521 \$153 \$8951 \$8912 \$8723 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31522 \$16 \$7378 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31523 \$16 \$7521 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31524 \$153 \$8782 \$8885 \$8604 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31525 \$16 \$8715 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31526 \$153 \$8997 \$8535 \$8715 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31528 \$16 \$8828 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31529 \$16 \$7521 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31530 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$31531 \$153 \$8897 \$8912 \$8604 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31532 \$153 \$8897 \$8535 \$8950 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31533 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$31534 \$16 \$8715 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31535 \$153 \$8857 \$8668 \$8715 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31536 \$16 \$8950 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31539 \$153 \$8911 \$8668 \$8950 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31540 \$153 \$8857 \$8638 \$8565 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31541 \$16 \$8950 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31542 \$153 \$8911 \$8912 \$8565 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31543 \$153 \$8952 \$8668 \$8828 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31545 \$16 \$7154 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31547 \$153 \$8913 \$8642 \$8950 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31548 \$16 \$8828 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31549 \$16 \$6909 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31550 \$16 \$8117 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31551 \$153 \$8914 \$8642 \$9026 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31552 \$153 \$8952 \$8885 \$8565 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31554 \$16 \$8950 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31555 \$153 \$8913 \$8912 \$8513 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31556 \$16 \$9026 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31557 \$153 \$8930 \$8642 \$8828 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31558 \$16 \$8025 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31559 \$16 \$7502 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31560 \$16 \$8118 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31562 \$153 \$8930 \$8885 \$8513 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31563 \$16 \$8828 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31564 \$16 \$8436 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31565 \$16 \$8715 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31566 \$153 \$8953 \$8669 \$8715 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31567 \$16 \$8365 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31569 \$153 \$8914 \$8726 \$8513 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31570 \$16 \$8828 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31571 \$153 \$8829 \$8669 \$8828 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31572 \$153 \$8953 \$8638 \$8515 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31573 \$16 \$7226 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31574 \$16 \$6935 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31575 \$16 \$8169 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31576 \$16 \$7000 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31578 \$16 \$8436 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31579 \$16 \$8436 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31580 \$16 \$8828 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31581 \$16 \$8715 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31582 \$153 \$8830 \$8740 \$8828 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31583 \$153 \$8858 \$8740 \$8715 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31584 \$16 \$8177 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31585 \$153 \$8831 \$8740 \$9026 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31587 \$16 \$6915 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31588 \$16 \$6910 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31590 \$153 \$8858 \$8638 \$8567 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31591 \$16 \$9026 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31592 \$16 \$7212 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31593 \$16 \$6910 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31594 \$153 \$8832 \$8740 \$8950 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31595 \$153 \$153 \$8726 \$8981 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31597 \$16 \$8635 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31598 \$16 \$8516 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31599 \$16 \$8950 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31600 \$153 \$8859 \$8740 \$8724 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31602 \$16 \$8670 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31603 \$153 \$9747 \$7041 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$31604 \$153 \$8859 \$8457 \$8567 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31605 \$16 \$9747 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31606 \$16 \$8671 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31607 \$16 \$6732 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31608 \$16 \$8568 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31610 \$16 \$8890 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31612 \$16 \$8724 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31614 \$153 \$8983 \$8744 \$8890 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31616 \$153 \$8915 \$8744 \$8886 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31619 \$153 \$8983 \$8277 \$8569 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31620 \$153 \$8817 \$8804 \$8569 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31622 \$153 \$8915 \$8727 \$8569 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31623 \$153 \$8984 \$8727 \$9097 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31624 \$16 \$8890 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31625 \$16 \$8886 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31627 \$153 \$8833 \$8743 \$8686 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31628 \$153 \$8986 \$8743 \$8728 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31630 \$153 \$8985 \$8789 \$9097 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31631 \$153 \$8860 \$8789 \$8569 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31632 \$16 \$8728 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31633 \$16 \$8686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31635 \$16 \$8728 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31636 \$153 \$8954 \$8586 \$8816 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31637 \$16 \$6987 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31638 \$16 \$6987 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31639 \$153 \$8684 \$8586 \$8898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31641 \$153 \$8742 \$8586 \$8886 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31642 \$153 \$8899 \$8277 \$8887 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31643 \$16 \$8898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31645 \$153 \$8987 \$8610 \$8887 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31646 \$16 \$8890 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31647 \$153 \$8888 \$8727 \$8424 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31648 \$16 \$8886 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31649 \$16 \$8635 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31651 \$153 \$8931 \$8587 \$8816 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31653 \$153 \$9003 \$8587 \$8890 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31654 \$16 \$8816 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31655 \$16 \$8890 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31656 \$153 \$8931 \$8804 \$8685 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31657 \$16 \$7071 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31658 \$153 \$8889 \$8609 \$8898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31661 \$153 \$8802 \$8609 \$8890 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31662 \$16 \$8898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31663 \$153 \$8888 \$8609 \$8886 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31664 \$16 \$8890 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31665 \$153 \$8803 \$8609 \$8816 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31667 \$153 \$8889 \$8789 \$8424 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31668 \$16 \$7502 \$8357 \$9004 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$31669 \$16 \$8816 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31671 \$16 \$8886 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31672 \$153 \$9005 \$8464 \$8890 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31673 \$16 \$7502 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31674 \$153 \$8932 \$8464 \$8898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31676 \$16 \$8890 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31677 \$16 \$8898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31679 \$153 \$9006 \$8464 \$8816 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31680 \$153 \$8805 \$8464 \$8886 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31681 \$16 \$8816 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31683 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$31684 \$16 \$8556 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31685 \$16 \$8886 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31687 \$153 \$9007 \$8611 \$8890 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31689 \$153 \$8933 \$8611 \$8816 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31690 \$153 \$8933 \$8804 \$8572 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31691 \$16 \$8816 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31693 \$153 \$8835 \$8611 \$8898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31694 \$16 \$8890 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31697 \$153 \$8834 \$8611 \$8886 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31698 \$16 \$8898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31699 \$16 \$8886 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31700 \$153 \$8750 \$8612 \$8890 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31701 \$153 \$8988 \$8612 \$8816 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31703 \$16 \$8890 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31704 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$31705 \$153 \$8988 \$8804 \$8613 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31707 \$153 \$8934 \$8612 \$8898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31708 \$16 \$8816 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31709 \$16 \$8728 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31710 \$16 \$8686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31711 \$153 \$8934 \$8789 \$8613 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31712 \$16 \$8898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31713 \$153 \$8836 \$8557 \$8886 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31715 \$153 \$9008 \$8818 \$8989 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31717 \$153 \$8970 \$8610 \$8989 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31719 \$153 \$8790 \$8804 \$8688 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31721 \$153 \$9011 \$8557 \$8890 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31723 \$16 \$8890 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31724 \$16 \$8898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31726 \$153 \$8837 \$8557 \$8898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31727 \$153 \$8957 \$8340 \$7065 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31728 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31729 \$153 \$8788 \$8340 \$7366 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31730 \$16 \$10143 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31731 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31734 \$153 \$8955 \$8340 \$7066 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31735 \$153 \$10143 \$7239 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$31736 \$153 \$8956 \$8340 \$6582 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31737 \$16 \$7129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31740 \$16 \$8839 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31741 \$16 \$10135 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31742 \$153 \$10135 \$7328 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$31743 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31745 \$16 \$8936 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31746 \$153 \$8990 \$9174 \$8126 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31747 \$153 \$8991 \$8676 \$8958 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31748 \$153 \$8618 \$7065 \$8538 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31751 \$153 \$8959 \$8935 \$8936 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31752 \$153 \$8935 \$7484 \$8791 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$31753 \$153 \$8991 \$8935 \$8807 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31754 \$16 \$8807 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31755 \$16 \$7067 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31756 \$16 \$7344 \$16 \$153 \$8958 VNB sky130_fd_sc_hd__inv_1
X$31759 \$16 \$7328 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31760 \$16 \$8719 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31761 \$16 \$8673 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31763 \$16 \$8820 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31764 \$16 \$7082 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31765 \$16 \$7350 \$8819 \$8971 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$31766 \$153 \$8861 \$6582 \$8373 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31767 \$153 \$8900 \$7551 \$8971 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$31768 \$16 \$8936 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31770 \$153 \$8862 \$8900 \$8807 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31773 \$16 \$9031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31775 \$16 \$8936 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31776 \$153 \$9012 \$8842 \$8891 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31777 \$153 \$8862 \$8676 \$8891 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31779 \$153 \$9013 \$8972 \$8936 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31780 \$153 \$8916 \$8917 \$9324 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31781 \$16 \$8821 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31783 \$153 \$8620 \$3916 \$8558 \$8863 \$8808 \$8560 \$8593 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$31784 \$153 \$8841 \$8972 \$8807 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31785 \$153 \$9013 \$8842 \$8840 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31786 \$16 \$8863 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31788 \$153 \$8972 \$8794 \$8918 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$31790 \$153 \$8937 \$8869 \$8992 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$31791 \$153 \$8919 \$9174 \$7994 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31792 \$153 \$9014 \$8937 \$8936 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31793 \$153 \$8901 \$8676 \$8843 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31795 \$16 \$7130 \$8819 \$8992 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$31796 \$153 \$8901 \$8937 \$8807 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31798 \$153 \$8938 \$8621 \$7082 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31800 \$153 \$8938 \$7065 \$8525 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31801 \$153 \$8793 \$7490 \$8525 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31803 \$153 \$9015 \$9047 \$8993 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31804 \$153 \$8864 \$8621 \$7067 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31806 \$16 \$7489 \$8960 \$8973 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$31807 \$153 \$9050 \$7686 \$8973 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$31808 \$153 \$8864 \$6582 \$8525 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31810 \$153 \$8865 \$8677 \$7239 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31811 \$153 \$8961 \$8677 \$7067 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31812 \$153 \$8865 \$7482 \$8574 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31813 \$153 \$8961 \$6582 \$8574 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31814 \$153 \$8866 \$8677 \$7387 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31815 \$16 \$8936 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31817 \$153 \$8809 \$8677 \$7082 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31818 \$153 \$8866 \$7490 \$8574 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31819 \$16 \$7082 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31820 \$16 \$7429 \$8960 \$8974 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$31821 \$16 \$8808 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31822 \$16 \$7429 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31823 \$153 \$9053 \$7614 \$8974 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$31824 \$16 \$7082 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31826 \$153 \$8867 \$8733 \$7082 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31827 \$16 \$7614 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31828 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$31829 \$153 \$8867 \$7065 \$8691 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31830 \$16 \$8807 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31831 \$153 \$8770 \$7215 \$8691 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31832 \$16 \$7067 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31833 \$16 \$8936 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31836 \$153 \$8962 \$9053 \$8936 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31837 \$16 \$7429 \$16 \$153 \$8920 VNB sky130_fd_sc_hd__inv_1
X$31838 \$153 \$8921 \$8733 \$7067 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31839 \$16 \$8265 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31840 \$153 \$8921 \$6582 \$8691 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31841 \$16 \$7429 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31843 \$16 \$8704 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31844 \$16 \$7239 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31846 \$16 \$7498 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31847 \$153 \$8868 \$8733 \$7239 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31848 \$16 \$7267 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31849 \$16 \$9188 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31851 \$16 \$7498 \$8960 \$8975 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$31852 \$153 \$9054 \$7267 \$8975 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$31853 \$153 \$8868 \$7482 \$8691 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31854 \$16 \$8734 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31856 \$16 \$8936 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31857 \$16 \$10383 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31859 \$153 \$9017 \$9054 \$8936 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31860 \$16 \$7607 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31861 \$16 \$8735 \$8473 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$31862 \$16 \$8822 \$7484 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$31863 \$16 \$8822 \$7903 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$31864 \$16 \$8902 \$16 \$153 \$8822 VNB sky130_fd_sc_hd__clkbuf_2
X$31866 \$153 \$8994 \$8676 \$9151 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31867 \$16 \$8340 \$16 \$153 \$8902 VNB sky130_fd_sc_hd__clkbuf_2
X$31868 \$16 \$8902 \$16 \$153 \$8735 VNB sky130_fd_sc_hd__clkbuf_2
X$31869 \$16 \$8823 \$7267 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$31870 \$16 \$8902 \$16 \$153 \$9055 VNB sky130_fd_sc_hd__clkbuf_2
X$31872 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31873 \$16 \$8902 \$16 \$153 \$8823 VNB sky130_fd_sc_hd__clkbuf_2
X$31874 \$153 \$8904 \$8869 \$8903 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$31875 \$16 \$7130 \$8824 \$8903 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$31876 \$16 \$8416 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31877 \$153 \$9018 \$8904 \$8927 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31878 \$153 \$8939 \$8904 \$8893 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31880 \$16 \$8927 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31881 \$153 \$8939 \$8996 \$8892 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31883 \$16 \$7130 \$16 \$153 \$8892 VNB sky130_fd_sc_hd__inv_1
X$31884 \$16 \$8893 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31885 \$153 \$8922 \$7484 \$8870 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$31886 \$16 \$9035 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31887 \$16 \$7375 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31888 \$16 \$8719 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31889 \$153 \$8905 \$8904 \$8844 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31890 \$16 \$8187 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31891 \$16 \$8673 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31893 \$16 \$8673 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31894 \$153 \$8905 \$8965 \$8892 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31895 \$16 \$8844 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31897 \$16 \$8820 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31898 \$16 \$8927 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31899 \$153 \$8940 \$8922 \$8844 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31900 \$153 \$9020 \$8922 \$8927 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31901 \$16 \$7344 \$16 \$153 \$8906 VNB sky130_fd_sc_hd__inv_1
X$31903 \$153 \$8940 \$8965 \$8906 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31905 \$153 \$8811 \$8922 \$8893 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31906 \$16 \$9150 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31907 \$16 \$7668 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31908 \$16 \$7495 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31909 \$16 \$8893 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31910 \$153 \$8976 \$8977 \$8906 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31911 \$153 \$8872 \$8923 \$8906 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31912 \$16 \$8844 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31914 \$153 \$8941 \$8812 \$8844 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31916 \$153 \$8963 \$8812 \$8927 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31917 \$16 \$7495 \$8824 \$8873 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$31918 \$153 \$8941 \$8965 \$8995 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31919 \$153 \$8942 \$8812 \$8879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31920 \$16 \$8220 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31923 \$16 \$8844 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31924 \$153 \$8942 \$8923 \$8995 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31925 \$16 \$8879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31927 \$153 \$8924 \$8874 \$8879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31928 \$153 \$9036 \$8874 \$8844 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31930 \$16 \$7495 \$16 \$153 \$8943 VNB sky130_fd_sc_hd__inv_1
X$31931 \$16 \$7495 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31932 \$16 \$8291 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31933 \$16 \$8879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31935 \$16 \$8893 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31936 \$16 \$8927 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31937 \$153 \$8964 \$8874 \$8927 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31938 \$153 \$8925 \$8874 \$8893 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31939 \$153 \$8926 \$7686 \$8875 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$31940 \$16 \$7686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31942 \$16 \$8879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31944 \$153 \$8925 \$8996 \$8943 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31945 \$153 \$8944 \$8926 \$8844 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31946 \$153 \$8847 \$8926 \$8879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31948 \$153 \$8944 \$8965 \$8846 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31949 \$16 \$8879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31951 \$153 \$8908 \$8772 \$8907 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$31952 \$16 \$7952 \$8825 \$8907 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$31954 \$153 \$8850 \$8908 \$8927 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31955 \$153 \$8814 \$8908 \$8879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31957 \$16 \$8927 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31959 \$16 \$8844 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31960 \$16 \$8893 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31961 \$153 \$8945 \$8908 \$8844 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31962 \$153 \$8966 \$8908 \$8893 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31963 \$153 \$8945 \$8965 \$8849 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31964 \$16 \$8291 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31965 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$31966 \$16 \$7429 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31968 \$16 \$7429 \$8825 \$8876 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$31969 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$31970 \$16 \$8927 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31971 \$16 \$8844 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31972 \$153 \$9022 \$8877 \$8927 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31973 \$153 \$8946 \$8877 \$8844 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31974 \$16 \$7431 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31975 \$16 \$7429 \$16 \$153 \$8852 VNB sky130_fd_sc_hd__inv_1
X$31976 \$16 \$7267 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31977 \$16 \$8893 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31979 \$16 \$8879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31981 \$153 \$8880 \$8877 \$8879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31982 \$153 \$9023 \$8877 \$8893 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31983 \$153 \$8880 \$8923 \$8852 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31984 \$153 \$8929 \$7267 \$8928 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$31985 \$16 \$8879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31987 \$16 \$7498 \$8825 \$8928 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$31988 \$153 \$8967 \$8929 \$8893 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31989 \$153 \$8894 \$8929 \$8879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31990 \$153 \$8967 \$8996 \$8947 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31991 \$153 \$8894 \$8923 \$8947 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$31994 \$16 \$8428 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31995 \$16 \$7498 \$16 \$153 \$8947 VNB sky130_fd_sc_hd__inv_1
X$31996 \$16 \$9154 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$31998 \$153 \$8968 \$8929 \$9154 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$31999 \$153 \$8853 \$8929 \$8844 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32000 \$153 \$8968 \$9103 \$8947 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32001 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$32003 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$32004 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$32006 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$32007 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$32008 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$32009 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$32010 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$32011 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$32012 \$153 \$8978 \$8895 \$8950 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32013 \$153 \$9037 \$8895 \$8715 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32014 \$16 \$8950 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32015 \$16 \$8715 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32016 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$32017 \$16 \$6915 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32018 \$153 \$9061 \$8737 \$9025 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32021 \$153 \$9104 \$8895 \$8828 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32022 \$153 \$9037 \$8638 \$8882 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32023 \$153 \$9062 \$8638 \$8679 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32024 \$153 \$9104 \$8885 \$8882 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32025 \$16 \$8828 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32026 \$153 \$9105 \$8895 \$8436 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32027 \$16 \$7545 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32029 \$16 \$7545 \$16 \$153 \$9025 VNB sky130_fd_sc_hd__inv_1
X$32030 \$153 \$9063 \$8457 \$8882 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32031 \$153 \$9064 \$8726 \$8679 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32032 \$153 \$9105 \$8209 \$8882 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32033 \$153 \$9065 \$8209 \$8679 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32034 \$16 \$7545 \$8577 \$9157 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$32037 \$153 \$9196 \$7333 \$9067 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$32038 \$16 \$7237 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32039 \$16 \$7545 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32040 \$153 \$9066 \$8722 \$9026 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32041 \$16 \$6988 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32043 \$153 \$9106 \$9196 \$9129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32044 \$16 \$7378 \$8577 \$9067 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$32047 \$16 \$9026 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32048 \$153 \$9038 \$8726 \$8883 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32049 \$16 \$7378 \$16 \$153 \$8883 VNB sky130_fd_sc_hd__inv_1
X$32050 \$16 \$9129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32052 \$153 \$8951 \$8533 \$8950 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32053 \$153 \$8717 \$8533 \$9026 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32054 \$153 \$9106 \$8737 \$8883 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32057 \$16 \$9026 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32059 \$16 \$8828 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32060 \$153 \$9135 \$8885 \$9136 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32061 \$16 \$8950 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32063 \$153 \$9068 \$8535 \$9026 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32065 \$153 \$9158 \$9130 \$8436 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32068 \$16 \$9026 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32069 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$32070 \$16 \$8436 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32073 \$16 \$6909 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32074 \$153 \$8997 \$8638 \$8604 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32075 \$16 \$8715 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32076 \$153 \$9107 \$9131 \$8715 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32077 \$153 \$9068 \$8726 \$8604 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32078 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$32080 \$153 \$9069 \$8737 \$9027 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32082 \$153 \$9107 \$8638 \$9027 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32083 \$16 \$7071 \$8504 \$9028 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$32084 \$16 \$7071 \$16 \$153 \$9027 VNB sky130_fd_sc_hd__inv_1
X$32085 \$16 \$7071 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32086 \$153 \$9131 \$7154 \$9028 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$32087 \$16 \$7071 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32089 \$153 \$9130 \$7156 \$9070 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$32091 \$16 \$6909 \$8504 \$9070 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$32092 \$16 \$9220 \$16 \$153 \$8504 VNB sky130_fd_sc_hd__clkbuf_2
X$32093 \$16 \$8715 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32094 \$153 \$8998 \$9039 \$8715 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32095 \$153 \$9071 \$9039 \$9026 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32096 \$16 \$9026 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32097 \$153 \$9071 \$8726 \$9029 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32098 \$16 \$7973 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32101 \$153 \$9108 \$9039 \$8580 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32102 \$16 \$8118 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32104 \$16 \$7502 \$8504 \$9040 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$32105 \$153 \$9039 \$8365 \$9040 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$32106 \$153 \$9108 \$8194 \$9029 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32107 \$16 \$7502 \$16 \$153 \$9029 VNB sky130_fd_sc_hd__inv_1
X$32108 \$16 \$8580 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32110 \$153 \$9137 \$8737 \$9029 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32111 \$153 \$8999 \$8669 \$8950 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32113 \$16 \$8724 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32114 \$153 \$8800 \$8669 \$9026 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32115 \$153 \$8999 \$8912 \$8515 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32116 \$16 \$8950 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32119 \$16 \$9026 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32120 \$153 \$9109 \$9160 \$9026 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32122 \$153 \$9000 \$9160 \$8436 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32123 \$153 \$9109 \$8726 \$9072 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32124 \$153 \$9000 \$8209 \$9072 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32125 \$16 \$7072 \$8504 \$9073 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$32127 \$153 \$9160 \$7165 \$9073 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$32128 \$153 \$153 \$8885 \$8981 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32129 \$153 \$153 \$8638 \$8981 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32130 \$153 \$153 \$8194 \$8981 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32131 \$16 \$16 \$153 VNB sky130_fd_sc_hd__conb_1
X$32133 \$16 \$8950 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32134 \$16 \$7288 \$16 \$153 \$8981 VNB sky130_fd_sc_hd__clkbuf_2
X$32136 \$16 \$7124 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32137 \$153 \$153 \$8912 \$8981 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32139 \$16 \$7288 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32140 \$16 \$6988 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32141 \$16 \$6888 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32142 \$153 \$9138 \$6784 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$32143 \$16 \$6719 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32145 \$153 \$8672 \$8743 \$8890 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32146 \$153 \$8984 \$8743 \$8886 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32148 \$153 \$9074 \$8743 \$8816 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32149 \$16 \$9138 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32150 \$16 \$8816 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32151 \$153 \$9074 \$8804 \$9097 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32152 \$153 \$9096 \$8743 \$8647 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32153 \$16 \$8886 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32157 \$153 \$9096 \$8614 \$9097 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32158 \$16 \$8647 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32159 \$153 \$8985 \$8743 \$8898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32160 \$16 \$6915 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32161 \$153 \$9110 \$8743 \$8556 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32162 \$16 \$8898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32163 \$16 \$7333 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32166 \$16 \$8556 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32167 \$16 \$8635 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32169 \$153 \$9139 \$8818 \$9185 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32170 \$16 \$7378 \$8635 \$9041 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$32171 \$153 \$9001 \$7333 \$9041 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$32172 \$153 \$9140 \$8818 \$9417 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32174 \$16 \$7378 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32175 \$16 \$7378 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32176 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$32177 \$16 \$7378 \$16 \$153 \$8887 VNB sky130_fd_sc_hd__inv_1
X$32178 \$16 \$8816 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32180 \$153 \$9110 \$8610 \$9097 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32181 \$153 \$8987 \$9001 \$8556 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32183 \$153 \$9163 \$9001 \$8686 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32184 \$153 \$8986 \$8818 \$9097 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32185 \$16 \$8556 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32186 \$16 \$8686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32188 \$153 \$9002 \$8587 \$8898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32190 \$153 \$9098 \$8587 \$8886 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32191 \$153 \$9002 \$8789 \$8685 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32193 \$153 \$9003 \$8277 \$8685 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32194 \$153 \$9098 \$8727 \$8685 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32197 \$16 \$8886 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32199 \$16 \$7071 \$16 \$153 \$9111 VNB sky130_fd_sc_hd__inv_1
X$32200 \$16 \$8898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32201 \$153 \$9141 \$8727 \$9111 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32202 \$16 \$7071 \$8357 \$9042 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$32203 \$153 \$9132 \$7154 \$9042 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$32204 \$153 \$9112 \$9132 \$8898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32207 \$16 \$8898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32208 \$153 \$9076 \$8365 \$9004 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$32209 \$153 \$9112 \$8789 \$9111 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32210 \$153 \$9142 \$8818 \$9111 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32211 \$16 \$8365 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32213 \$153 \$9005 \$8277 \$8687 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32214 \$16 \$9273 \$16 \$153 \$8357 VNB sky130_fd_sc_hd__clkbuf_2
X$32215 \$16 \$7502 \$16 \$153 \$9144 VNB sky130_fd_sc_hd__inv_1
X$32217 \$153 \$8932 \$8789 \$8687 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32218 \$153 \$9143 \$8789 \$9144 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32219 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$32220 \$16 \$7502 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32221 \$153 \$9113 \$9076 \$8686 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32222 \$153 \$9006 \$8804 \$8687 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32224 \$153 \$9113 \$8651 \$9144 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32226 \$16 \$8686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32227 \$16 \$7156 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32228 \$153 \$9077 \$7156 \$9043 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$32229 \$16 \$6909 \$8357 \$9043 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$32230 \$153 \$9007 \$8277 \$8572 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32231 \$153 \$9078 \$9077 \$8556 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32232 \$16 \$6909 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32233 \$16 \$6909 \$16 \$153 \$9146 VNB sky130_fd_sc_hd__inv_1
X$32236 \$16 \$7072 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32237 \$153 \$9145 \$8789 \$9146 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32238 \$16 \$8556 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32240 \$16 \$7072 \$8357 \$9030 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$32241 \$16 \$7165 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32243 \$153 \$9044 \$7165 \$9030 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$32244 \$153 \$9165 \$9077 \$8647 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32247 \$16 \$8647 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32248 \$153 \$9114 \$9077 \$8686 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32249 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$32250 \$153 \$9008 \$9044 \$8728 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32251 \$153 \$9114 \$8651 \$9146 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32252 \$153 \$9009 \$9044 \$8686 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32255 \$153 \$8970 \$9044 \$8556 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32256 \$153 \$9009 \$8651 \$8989 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32257 \$153 \$153 \$8610 \$9010 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32258 \$16 \$7072 \$16 \$153 \$8989 VNB sky130_fd_sc_hd__inv_1
X$32259 \$16 \$7288 \$16 \$153 \$9010 VNB sky130_fd_sc_hd__clkbuf_2
X$32260 \$153 \$153 \$8651 \$9010 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32262 \$153 \$153 \$8804 \$9010 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32263 \$16 \$16 \$153 VNB sky130_fd_sc_hd__conb_1
X$32264 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32265 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32267 \$153 \$9075 \$8340 \$7482 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32268 \$153 \$8657 \$9116 \$8807 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32269 \$153 \$9227 \$7067 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$32271 \$153 \$9011 \$8277 \$8688 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32272 \$16 \$8807 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32273 \$16 \$8936 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32274 \$153 \$9099 \$9116 \$8936 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32275 \$153 \$9079 \$9133 \$8126 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32277 \$16 \$7366 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32278 \$16 \$7327 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32280 \$153 \$8919 \$9116 \$9045 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32281 \$153 \$9147 \$9252 \$8126 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32282 \$16 \$9045 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32283 \$153 \$9116 \$7347 \$9166 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$32284 \$153 \$9046 \$9047 \$8126 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32286 \$16 \$7386 \$16 \$153 \$7994 VNB sky130_fd_sc_hd__inv_1
X$32288 \$153 \$9167 \$8935 \$9045 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32290 \$153 \$9080 \$8935 \$9214 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32291 \$153 \$9168 \$8935 \$9031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32292 \$16 \$7386 \$8819 \$9166 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$32293 \$16 \$9214 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32296 \$153 \$8959 \$8842 \$8958 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32297 \$16 \$8819 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32299 \$16 \$8819 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32300 \$153 \$9167 \$9174 \$8958 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32301 \$16 \$9045 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32302 \$153 \$9048 \$8900 \$9045 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32304 \$153 \$9012 \$8900 \$8936 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32306 \$153 \$9100 \$8900 \$9031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32307 \$153 \$9048 \$9174 \$8891 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32308 \$153 \$9100 \$9133 \$8891 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32310 \$153 \$9170 \$8972 \$9214 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32312 \$16 \$9045 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32315 \$153 \$9081 \$7668 \$9049 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$32316 \$153 \$9171 \$8972 \$9031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32317 \$153 \$9082 \$8972 \$9045 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32318 \$16 \$7667 \$8819 \$9049 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$32319 \$16 \$9045 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32321 \$153 \$9082 \$9174 \$8840 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32322 \$16 \$7495 \$8819 \$8918 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$32323 \$16 \$7495 \$16 \$153 \$8840 VNB sky130_fd_sc_hd__inv_1
X$32325 \$153 \$9101 \$8937 \$9045 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32326 \$153 \$9083 \$8937 \$9031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32327 \$153 \$9101 \$9174 \$8843 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32330 \$153 \$9014 \$8842 \$8843 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32331 \$16 \$9188 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32333 \$16 \$9031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32334 \$16 \$9031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32336 \$153 \$9117 \$9050 \$9031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32337 \$16 \$9214 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32338 \$153 \$9015 \$9050 \$9214 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32340 \$16 \$8936 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32341 \$153 \$9016 \$9050 \$8936 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32342 \$16 \$8794 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32343 \$16 \$7495 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32344 \$16 \$8807 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32345 \$153 \$9051 \$9050 \$8807 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32346 \$153 \$9016 \$8842 \$8993 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32347 \$153 \$9117 \$9133 \$8993 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32350 \$153 \$9051 \$8676 \$8993 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32351 \$153 \$9052 \$7693 \$9149 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$32352 \$16 \$7489 \$16 \$153 \$8993 VNB sky130_fd_sc_hd__inv_1
X$32354 \$153 \$9084 \$9052 \$9045 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32355 \$16 \$9045 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32356 \$16 \$9031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32357 \$16 \$7067 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32359 \$16 \$8807 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32361 \$153 \$9118 \$9052 \$8807 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32363 \$153 \$9085 \$9052 \$8936 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32365 \$153 \$9085 \$8842 \$9033 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32366 \$153 \$9032 \$9133 \$9033 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32368 \$16 \$7693 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32370 \$16 \$9214 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32372 \$16 \$9045 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32373 \$153 \$9175 \$9053 \$9214 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32374 \$153 \$9086 \$9053 \$9045 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32376 \$153 \$9086 \$9174 \$8920 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32377 \$153 \$9087 \$9053 \$8807 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32379 \$153 \$9175 \$9047 \$8920 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32380 \$153 \$8962 \$8842 \$8920 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32381 \$153 \$9087 \$8676 \$8920 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32382 \$16 \$9188 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32383 \$16 \$8344 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32384 \$16 \$9045 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32385 \$16 \$8498 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32386 \$153 \$9119 \$9054 \$9045 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32387 \$16 \$7306 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32388 \$16 \$7498 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32389 \$16 \$9214 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32391 \$153 \$9088 \$9054 \$9214 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32392 \$153 \$9088 \$9047 \$9151 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32393 \$16 \$7498 \$16 \$153 \$9151 VNB sky130_fd_sc_hd__inv_1
X$32394 \$153 \$9119 \$9174 \$9151 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32395 \$16 \$7462 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32396 \$16 \$8807 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32397 \$153 \$8994 \$9054 \$8807 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32398 \$16 \$9031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32400 \$153 \$9177 \$9054 \$9031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32401 \$153 \$9017 \$8842 \$9151 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32402 \$16 \$7130 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32403 \$16 \$9055 \$8627 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$32404 \$16 \$8869 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32405 \$16 \$9055 \$8250 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$32406 \$16 \$9055 \$7839 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$32407 \$153 \$9179 \$7347 \$9178 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$32408 \$16 \$9055 \$8820 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$32410 \$16 \$9055 \$8719 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$32411 \$16 \$9055 \$8731 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$32412 \$16 \$9134 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32413 \$153 \$9089 \$8904 \$9134 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32414 \$153 \$9120 \$9256 \$9152 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32415 \$153 \$9153 \$8923 \$9152 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32416 \$153 \$9019 \$8904 \$9035 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32418 \$16 \$9134 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32419 \$153 \$9018 \$9256 \$8892 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32420 \$153 \$9090 \$8904 \$9034 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32421 \$16 \$9055 \$9150 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$32422 \$16 \$7130 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32423 \$153 \$9056 \$8904 \$9154 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32425 \$153 \$9019 \$8977 \$8892 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32426 \$16 \$9154 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32427 \$16 \$9034 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32428 \$16 \$8313 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32429 \$153 \$9056 \$9103 \$8892 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32431 \$153 \$9121 \$8922 \$9034 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32432 \$153 \$8871 \$8923 \$8892 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32434 \$16 \$8844 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32436 \$153 \$9121 \$9059 \$8906 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32438 \$16 \$9035 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32439 \$153 \$8976 \$8922 \$9035 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32440 \$16 \$9034 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32441 \$16 \$7551 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32443 \$153 \$9123 \$9122 \$8995 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32444 \$16 \$7350 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32445 \$16 \$7996 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32446 \$16 \$8927 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32447 \$153 \$9124 \$9059 \$8995 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32448 \$16 \$9154 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32450 \$153 \$9102 \$8812 \$9154 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32451 \$153 \$9102 \$9103 \$8995 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32452 \$153 \$9125 \$8977 \$8995 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32454 \$16 \$7667 \$16 \$153 \$8995 VNB sky130_fd_sc_hd__inv_1
X$32456 \$153 \$9021 \$8812 \$8893 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32457 \$16 \$9134 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32458 \$16 \$8794 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32459 \$16 \$9034 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32461 \$153 \$9124 \$8812 \$9034 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32462 \$153 \$9021 \$8996 \$8995 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32463 \$16 \$9035 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32465 \$153 \$9036 \$8965 \$8943 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32466 \$153 \$9057 \$8874 \$9035 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32468 \$16 \$7667 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32469 \$16 \$8266 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32470 \$153 \$9057 \$8977 \$8943 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32471 \$16 \$9134 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32472 \$16 \$9154 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32473 \$153 \$9181 \$8874 \$9154 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32474 \$153 \$8924 \$8923 \$8943 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32475 \$153 \$8964 \$9256 \$8943 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32479 \$16 \$8291 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32481 \$16 \$7489 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32482 \$16 \$8893 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32483 \$16 \$7489 \$16 \$153 \$8846 VNB sky130_fd_sc_hd__inv_1
X$32484 \$16 \$9035 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32485 \$153 \$9182 \$8926 \$9035 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32486 \$153 \$9091 \$8926 \$8893 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32487 \$153 \$9155 \$9122 \$8943 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32488 \$16 \$8032 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32491 \$16 \$8772 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32492 \$153 \$9058 \$9103 \$8846 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32493 \$16 \$7952 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32495 \$16 \$9034 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32496 \$153 \$9092 \$8908 \$9034 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32497 \$153 \$9091 \$8996 \$8846 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32499 \$153 \$9092 \$9059 \$8849 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32500 \$16 \$7540 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32503 \$16 \$7952 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32504 \$16 \$7952 \$16 \$153 \$8849 VNB sky130_fd_sc_hd__inv_1
X$32505 \$16 \$9134 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32506 \$153 \$9093 \$9103 \$8849 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32507 \$16 \$9035 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32508 \$153 \$9126 \$8908 \$9035 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32509 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$32511 \$153 \$8966 \$8996 \$8849 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32512 \$153 \$9126 \$8977 \$8849 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32514 \$153 \$9094 \$9122 \$8849 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32515 \$16 \$9154 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32516 \$153 \$9183 \$8877 \$9154 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32517 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$32518 \$153 \$9022 \$9256 \$8852 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32519 \$16 \$7431 \$8825 \$9156 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$32520 \$153 \$8946 \$8965 \$8852 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32521 \$16 \$9035 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32524 \$153 \$9127 \$8877 \$9035 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32525 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$32526 \$153 \$9060 \$9059 \$8852 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32527 \$153 \$9023 \$8996 \$8852 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32528 \$153 \$9127 \$8977 \$8852 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32529 \$16 \$8927 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32530 \$16 \$8893 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32531 \$16 \$8927 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32535 \$153 \$9024 \$8929 \$8927 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32536 \$153 \$9128 \$8929 \$9134 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32537 \$153 \$9024 \$9256 \$8947 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32538 \$153 \$9128 \$9122 \$8947 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32539 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$32542 \$16 \$9034 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32544 \$153 \$9184 \$8929 \$9034 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32545 \$16 \$9035 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32546 \$153 \$9095 \$8929 \$9035 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32548 \$153 \$9095 \$8977 \$8947 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32549 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$32552 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$32553 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$32555 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$32556 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$32557 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$32558 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$32559 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$32560 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$32561 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$32562 \$153 \$678 \$511 \$17 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32563 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$32565 \$153 \$709 \$234 \$598 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32567 \$153 \$967 \$234 \$763 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32568 \$153 \$709 \$511 \$263 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32569 \$153 \$678 \$102 \$598 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32570 \$153 \$617 \$30 \$598 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32572 \$153 \$511 \$753 \$780 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$32573 \$16 \$263 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32576 \$153 \$679 \$511 \$419 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32577 \$153 \$530 \$394 \$598 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32578 \$153 \$679 \$349 \$598 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32579 \$153 \$618 \$59 \$598 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32580 \$16 \$710 \$16 \$153 \$598 VNB sky130_fd_sc_hd__inv_1
X$32582 \$16 \$419 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32583 \$153 \$680 \$661 \$419 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32585 \$153 \$711 \$661 \$263 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32586 \$153 \$680 \$349 \$649 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32587 \$153 \$764 \$394 \$649 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32588 \$16 \$419 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32589 \$16 \$263 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32590 \$16 \$783 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32591 \$16 \$710 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32593 \$16 \$249 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32594 \$16 \$783 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32595 \$153 \$661 \$662 \$599 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$32596 \$153 \$726 \$102 \$649 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32597 \$153 \$711 \$234 \$649 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32598 \$16 \$662 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32600 \$16 \$582 \$537 \$619 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$32601 \$16 \$754 \$16 \$153 \$649 VNB sky130_fd_sc_hd__inv_1
X$32602 \$153 \$663 \$561 \$783 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32603 \$16 \$754 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32604 \$16 \$503 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32607 \$153 \$712 \$59 \$903 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32608 \$153 \$66 \$541 \$533 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$32609 \$153 \$714 \$755 \$17 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32610 \$153 \$317 \$349 \$96 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32611 \$153 \$712 \$755 \$184 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32613 \$16 \$17 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32614 \$16 \$58 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32615 \$153 \$453 \$377 \$96 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32617 \$153 \$67 \$454 \$621 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$32618 \$153 \$620 \$561 \$96 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32619 \$16 \$184 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32621 \$16 \$504 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32622 \$16 \$395 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32624 \$153 \$785 \$817 \$419 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32625 \$153 \$681 \$561 \$639 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32626 \$153 \$68 \$1525 \$622 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$32627 \$16 \$419 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32629 \$16 \$503 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32630 \$16 \$1525 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32631 \$153 \$786 \$664 \$249 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32632 \$16 \$419 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32635 \$153 \$682 \$664 \$184 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32636 \$153 \$682 \$59 \$765 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32637 \$16 \$184 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32639 \$153 \$683 \$664 \$17 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32640 \$16 \$249 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32641 \$16 \$58 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32642 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$32644 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$32645 \$153 \$683 \$102 \$765 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32646 \$153 \$564 \$664 \$419 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32647 \$16 \$1551 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32648 \$153 \$650 \$756 \$58 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32649 \$16 \$419 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32650 \$16 \$356 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32653 \$153 \$190 \$684 \$623 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$32654 \$16 \$58 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32655 \$16 \$537 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32657 \$16 \$691 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32658 \$153 \$727 \$756 \$17 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32659 \$153 \$650 \$30 \$651 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32660 \$16 \$684 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32661 \$16 \$17 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32662 \$16 \$1508 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32664 \$16 \$504 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32666 \$153 \$727 \$102 \$651 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32667 \$16 \$419 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32668 \$153 \$640 \$583 \$17 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32669 \$16 \$849 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32671 \$16 \$715 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32672 \$16 \$17 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32673 \$153 \$536 \$349 \$766 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32674 \$153 \$640 \$102 \$766 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32675 \$153 \$624 \$377 \$766 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32677 \$16 \$249 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32679 \$153 \$728 \$583 \$184 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32680 \$153 \$381 \$234 \$172 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32681 \$153 \$728 \$59 \$766 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32682 \$153 \$625 \$30 \$766 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32683 \$16 \$652 \$16 \$153 \$766 VNB sky130_fd_sc_hd__inv_1
X$32685 \$16 \$184 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32687 \$153 \$71 \$757 \$789 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$32688 \$16 \$685 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32689 \$153 \$686 \$506 \$419 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32690 \$16 \$716 \$715 \$729 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$32692 \$16 \$419 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32693 \$153 \$686 \$349 \$432 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32694 \$16 \$652 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32695 \$16 \$715 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32696 \$16 \$184 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32698 \$153 \$516 \$506 \$184 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32699 \$153 \$730 \$561 \$432 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32700 \$16 \$716 \$16 \$153 \$432 VNB sky130_fd_sc_hd__inv_1
X$32702 \$153 \$586 \$454 \$790 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$32703 \$16 \$454 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32704 \$16 \$585 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32705 \$153 \$626 \$35 \$641 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32707 \$153 \$687 \$586 \$209 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32708 \$153 \$731 \$586 \$187 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32709 \$153 \$687 \$346 \$641 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32710 \$153 \$731 \$54 \$641 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32711 \$16 \$209 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32712 \$16 \$280 \$16 \$153 \$641 VNB sky130_fd_sc_hd__inv_1
X$32714 \$16 \$280 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32715 \$153 \$717 \$586 \$358 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32717 \$153 \$717 \$253 \$641 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32718 \$153 \$718 \$586 \$18 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32719 \$16 \$358 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32721 \$153 \$688 \$586 \$60 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32723 \$16 \$18 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32724 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$32725 \$153 \$518 \$586 \$212 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32726 \$153 \$688 \$104 \$641 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32728 \$153 \$732 \$758 \$358 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32729 \$16 \$60 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32730 \$16 \$212 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32734 \$16 \$754 \$16 \$153 \$175 VNB sky130_fd_sc_hd__inv_1
X$32735 \$153 \$732 \$253 \$767 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32737 \$16 \$358 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32738 \$153 \$185 \$430 \$665 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$32739 \$153 \$519 \$185 \$358 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32740 \$16 \$582 \$507 \$665 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$32743 \$153 \$570 \$253 \$175 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32744 \$153 \$540 \$54 \$105 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32746 \$153 \$719 \$587 \$18 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32749 \$16 \$293 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32750 \$153 \$653 \$587 \$187 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32751 \$16 \$710 \$16 \$153 \$600 VNB sky130_fd_sc_hd__inv_1
X$32752 \$16 \$18 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32754 \$153 \$733 \$587 \$358 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32755 \$153 \$653 \$54 \$600 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32757 \$16 \$187 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32758 \$16 \$358 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32759 \$16 \$555 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32761 \$153 \$689 \$587 \$60 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32762 \$153 \$734 \$587 \$209 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32763 \$153 \$689 \$104 \$600 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32764 \$16 \$356 \$555 \$601 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$32765 \$16 \$60 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32768 \$16 \$209 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32769 \$16 \$555 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32770 \$16 \$535 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32771 \$16 \$507 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32772 \$16 \$356 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32773 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$32775 \$153 \$735 \$690 \$18 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32776 \$153 \$654 \$690 \$358 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32777 \$16 \$18 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32778 \$153 \$654 \$253 \$655 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32779 \$16 \$18 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32782 \$16 \$358 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32783 \$16 \$691 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32785 \$16 \$351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32786 \$16 \$1264 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32787 \$153 \$642 \$690 \$60 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32788 \$16 \$1048 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32789 \$153 \$736 \$690 \$73 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32792 \$153 \$736 \$215 \$655 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32793 \$153 \$642 \$104 \$655 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32794 \$16 \$60 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32795 \$153 \$877 \$347 \$655 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32796 \$153 \$720 \$521 \$187 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32797 \$153 \$627 \$347 \$769 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32798 \$16 \$187 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32800 \$16 \$899 \$16 \$153 \$769 VNB sky130_fd_sc_hd__inv_1
X$32801 \$16 \$899 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32802 \$153 \$792 \$521 \$358 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32804 \$153 \$692 \$521 \$73 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32805 \$16 \$358 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32806 \$16 \$73 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32807 \$153 \$692 \$215 \$769 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32808 \$16 \$716 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32810 \$16 \$588 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32813 \$16 \$757 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32814 \$16 \$685 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32815 \$153 \$421 \$757 \$666 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$32816 \$153 \$75 \$685 \$793 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$32817 \$153 \$522 \$421 \$73 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32818 \$16 \$588 \$946 \$666 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$32819 \$16 \$716 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32821 \$16 \$60 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32823 \$153 \$794 \$759 \$60 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32824 \$153 \$667 \$54 \$760 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32825 \$153 \$629 \$35 \$436 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32827 \$153 \$737 \$759 \$209 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32828 \$16 \$209 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32829 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$32831 \$153 \$602 \$421 \$358 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32832 \$153 \$737 \$346 \$760 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32833 \$153 \$770 \$347 \$760 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32834 \$16 \$358 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32835 \$16 \$273 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32836 \$153 \$693 \$422 \$273 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32837 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$32840 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$32841 \$16 \$241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32842 \$153 \$693 \$389 \$501 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32845 \$153 \$738 \$826 \$79 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32848 \$153 \$477 \$353 \$501 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32849 \$16 \$399 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32850 \$153 \$630 \$266 \$501 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32851 \$153 \$545 \$388 \$501 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32852 \$153 \$694 \$559 \$501 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32853 \$16 \$594 \$16 \$153 \$501 VNB sky130_fd_sc_hd__inv_1
X$32854 \$16 \$397 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32855 \$16 \$273 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32856 \$16 \$558 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32857 \$153 \$603 \$407 \$273 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32858 \$16 \$424 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32860 \$153 \$589 \$407 \$424 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32861 \$153 \$878 \$266 \$656 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32862 \$16 \$82 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32863 \$153 \$606 \$407 \$82 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32865 \$16 \$399 \$268 \$668 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$32867 \$153 \$669 \$389 \$657 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32868 \$16 \$273 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32869 \$153 \$407 \$595 \$668 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$32870 \$153 \$557 \$388 \$604 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32871 \$16 \$424 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32873 \$153 \$739 \$559 \$605 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32874 \$16 \$82 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32875 \$153 \$643 \$590 \$82 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32876 \$153 \$740 \$590 \$424 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32877 \$16 \$884 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32878 \$16 \$964 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32879 \$16 \$268 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32880 \$153 \$740 \$353 \$605 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32882 \$153 \$643 \$44 \$605 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32883 \$16 \$798 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32884 \$16 \$397 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32885 \$16 \$438 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32887 \$16 \$424 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32888 \$153 \$696 \$670 \$424 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32890 \$153 \$409 \$266 \$604 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32891 \$153 \$697 \$670 \$273 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32892 \$153 \$742 \$670 \$79 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32895 \$16 \$424 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32897 \$153 \$303 \$44 \$485 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32898 \$16 \$79 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32899 \$16 \$354 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32900 \$16 \$79 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32901 \$16 \$82 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32902 \$153 \$644 \$592 \$82 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32903 \$153 \$743 \$592 \$79 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32906 \$16 \$273 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32907 \$153 \$743 \$112 \$607 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32908 \$153 \$881 \$388 \$607 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32909 \$153 \$644 \$44 \$607 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32910 \$153 \$1000 \$266 \$607 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32911 \$16 \$306 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32913 \$153 \$698 \$21 \$607 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32914 \$16 \$306 \$268 \$487 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$32915 \$16 \$268 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32916 \$153 \$699 \$559 \$771 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32917 \$153 \$800 \$389 \$771 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32919 \$16 \$700 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32920 \$153 \$744 \$388 \$771 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32921 \$16 \$424 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32922 \$16 \$82 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32923 \$153 \$609 \$593 \$82 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32924 \$153 \$772 \$266 \$771 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32926 \$153 \$801 \$44 \$611 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32928 \$16 \$273 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32929 \$16 \$273 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32932 \$153 \$745 \$830 \$273 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32933 \$153 \$645 \$425 \$424 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32934 \$153 \$745 \$389 \$611 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32935 \$153 \$645 \$353 \$348 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32938 \$16 \$145 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32939 \$16 \$276 \$441 \$671 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$32942 \$153 \$425 \$723 \$802 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$32943 \$153 \$62 \$1600 \$671 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$32944 \$153 \$673 \$830 \$145 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32945 \$153 \$672 \$112 \$611 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32949 \$153 \$673 \$266 \$611 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32950 \$153 \$773 \$21 \$611 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32951 \$16 \$1600 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32952 \$16 \$594 \$369 \$632 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$32953 \$153 \$803 \$761 \$509 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32954 \$16 \$724 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32955 \$16 \$426 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32956 \$16 \$369 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32957 \$16 \$309 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32958 \$153 \$524 \$391 \$309 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32961 \$153 \$804 \$549 \$774 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32962 \$16 \$509 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32963 \$153 \$633 \$393 \$442 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32964 \$16 \$558 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32965 \$16 \$594 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32966 \$16 \$63 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32968 \$153 \$612 \$391 \$63 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32970 \$153 \$746 \$23 \$774 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32971 \$153 \$883 \$57 \$774 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32973 \$16 \$446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32974 \$153 \$701 \$596 \$446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32975 \$16 \$509 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32976 \$16 \$884 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32977 \$16 \$902 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32980 \$16 \$310 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32981 \$153 \$701 \$393 \$658 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32982 \$16 \$399 \$428 \$634 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$32983 \$153 \$702 \$596 \$310 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32985 \$153 \$560 \$398 \$658 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32986 \$153 \$747 \$23 \$658 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32987 \$153 \$307 \$549 \$258 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32988 \$16 \$309 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32989 \$153 \$748 \$762 \$309 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$32990 \$16 \$428 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32991 \$16 \$631 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32992 \$16 \$674 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32993 \$153 \$227 \$674 \$370 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$32995 \$153 \$339 \$703 \$258 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32996 \$16 \$149 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$32997 \$153 \$675 \$223 \$659 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$32998 \$16 \$798 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33001 \$153 \$704 \$427 \$309 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33002 \$153 \$704 \$703 \$502 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33003 \$16 \$446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33004 \$153 \$705 \$427 \$446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33005 \$16 \$63 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33006 \$16 \$258 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33007 \$16 \$149 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33009 \$153 \$705 \$393 \$502 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33010 \$16 \$509 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33011 \$16 \$310 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33012 \$153 \$707 \$706 \$149 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33013 \$153 \$749 \$706 \$310 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33014 \$16 \$310 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33015 \$153 \$749 \$223 \$775 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33017 \$153 \$660 \$57 \$502 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33019 \$153 \$750 \$676 \$309 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33021 \$153 \$646 \$676 \$310 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33022 \$16 \$309 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33023 \$16 \$446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33024 \$153 \$646 \$223 \$445 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33027 \$153 \$707 \$398 \$775 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33029 \$16 \$149 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33031 \$153 \$614 \$676 \$63 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33032 \$16 \$63 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33034 \$153 \$647 \$23 \$445 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33035 \$153 \$751 \$398 \$776 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33036 \$153 \$777 \$371 \$445 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33037 \$16 \$509 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33038 \$16 \$309 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33039 \$153 \$597 \$723 \$677 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$33041 \$153 \$778 \$703 \$779 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33042 \$16 \$276 \$615 \$635 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$33045 \$153 \$808 \$597 \$509 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33046 \$153 \$708 \$597 \$309 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33047 \$153 \$636 \$57 \$637 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33048 \$16 \$508 \$615 \$677 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$33049 \$16 \$508 \$16 \$153 \$637 VNB sky130_fd_sc_hd__inv_1
X$33050 \$153 \$708 \$703 \$637 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33052 \$16 \$509 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33053 \$153 \$616 \$597 \$149 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33054 \$16 \$178 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33056 \$16 \$446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33057 \$153 \$725 \$836 \$446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33059 \$16 \$310 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33060 \$153 \$648 \$597 \$310 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33062 \$153 \$752 \$836 \$310 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33063 \$153 \$648 \$223 \$637 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33064 \$153 \$752 \$223 \$779 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33065 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$33066 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$33069 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$33071 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$33072 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$33073 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$33074 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$33075 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$33076 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$33078 \$153 \$9061 \$9193 \$9129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33080 \$153 \$9284 \$9193 \$8950 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33081 \$16 \$9129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33082 \$153 \$9194 \$8194 \$9025 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33083 \$16 \$8950 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33086 \$153 \$9284 \$8912 \$9025 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33088 \$16 \$7381 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33089 \$16 \$8724 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33091 \$16 \$8724 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33092 \$153 \$9063 \$8895 \$8724 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33093 \$153 \$9195 \$9193 \$8724 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33095 \$153 \$9266 \$8726 \$9025 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33096 \$153 \$9195 \$8457 \$9025 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33097 \$153 \$9267 \$8209 \$9025 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33098 \$16 \$8436 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33099 \$153 \$9193 \$7237 \$9157 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$33100 \$153 \$9268 \$8912 \$8679 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33101 \$16 \$8715 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33103 \$153 \$8980 \$9196 \$8828 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33105 \$153 \$8909 \$9196 \$8436 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33106 \$153 \$9197 \$8638 \$8883 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33107 \$16 \$8436 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33108 \$153 \$9198 \$9196 \$8580 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33109 \$16 \$8828 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33110 \$16 \$7333 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33112 \$153 \$9368 \$8912 \$8883 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33113 \$16 \$8580 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33115 \$153 \$9198 \$8194 \$8883 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33116 \$153 \$9269 \$8457 \$9270 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33119 \$153 \$9219 \$8726 \$9136 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33120 \$153 \$9135 \$9130 \$8828 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33122 \$153 \$9286 \$9130 \$8724 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33123 \$153 \$9219 \$9130 \$9026 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33124 \$153 \$9199 \$9130 \$8580 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33125 \$16 \$9220 \$16 \$153 \$8577 VNB sky130_fd_sc_hd__clkbuf_2
X$33128 \$16 \$9026 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33129 \$153 \$9199 \$8194 \$9136 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33130 \$16 \$8580 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33131 \$16 \$8724 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33133 \$153 \$9287 \$9131 \$8436 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33134 \$16 \$6909 \$16 \$153 \$9136 VNB sky130_fd_sc_hd__inv_1
X$33135 \$153 \$9069 \$9131 \$9129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33136 \$16 \$9026 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33139 \$153 \$9271 \$8726 \$9027 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33140 \$16 \$8436 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33141 \$16 \$9129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33142 \$153 \$9221 \$9131 \$8950 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33143 \$153 \$9287 \$8209 \$9027 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33145 \$153 \$9221 \$8912 \$9027 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33146 \$16 \$8950 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33147 \$16 \$7973 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33148 \$16 \$7156 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33151 \$16 \$9220 \$16 \$153 \$9260 VNB sky130_fd_sc_hd__clkbuf_2
X$33152 \$16 \$9200 \$16 \$153 \$9220 VNB sky130_fd_sc_hd__clkbuf_2
X$33153 \$16 \$8580 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33154 \$16 \$9200 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33156 \$153 \$9243 \$9039 \$8828 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33157 \$153 \$9222 \$9039 \$8436 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33158 \$153 \$8998 \$8638 \$9029 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33159 \$16 \$8828 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33160 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$33162 \$153 \$9243 \$8885 \$9029 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33163 \$16 \$8436 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33164 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$33165 \$153 \$9222 \$8209 \$9029 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33166 \$16 \$7502 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33167 \$153 \$9137 \$9039 \$9129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33168 \$16 \$9026 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33170 \$16 \$9129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33171 \$153 \$9289 \$9039 \$8724 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33173 \$153 \$9159 \$9039 \$8950 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33174 \$153 \$9159 \$8912 \$9029 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33175 \$16 \$8950 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33177 \$16 \$8580 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33178 \$16 \$7992 \$16 \$153 \$9322 VNB sky130_fd_sc_hd__inv_1
X$33179 \$16 \$8715 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33180 \$153 \$9161 \$9160 \$8715 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33181 \$16 \$6753 \$9260 \$9290 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$33183 \$153 \$9244 \$9160 \$8580 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33184 \$16 \$7992 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33185 \$16 \$8177 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33186 \$153 \$9161 \$8638 \$9072 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33187 \$153 \$9244 \$8194 \$9072 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33188 \$16 \$9026 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33189 \$16 \$6753 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33190 \$16 \$7072 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33191 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$33193 \$16 \$7072 \$16 \$153 \$9072 VNB sky130_fd_sc_hd__inv_1
X$33194 \$153 \$9245 \$9160 \$8950 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33195 \$16 \$7165 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33196 \$16 \$7072 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33198 \$153 \$9223 \$9160 \$8724 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33199 \$153 \$9245 \$8912 \$9072 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33200 \$153 \$153 \$8209 \$8981 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33202 \$153 \$153 \$8737 \$8981 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33203 \$16 \$8724 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33204 \$16 \$7237 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33205 \$153 \$9202 \$7237 \$9201 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$33206 \$153 \$153 \$8457 \$8981 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33207 \$16 \$7545 \$8635 \$9201 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$33209 \$16 \$7545 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33210 \$16 \$8635 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33212 \$16 \$6794 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33213 \$153 \$9246 \$9202 \$8816 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33215 \$153 \$9224 \$9202 \$8890 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33217 \$153 \$9246 \$8804 \$9185 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33218 \$153 \$9203 \$8727 \$9185 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33219 \$16 \$7545 \$16 \$153 \$9185 VNB sky130_fd_sc_hd__inv_1
X$33220 \$16 \$8890 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33222 \$16 \$6988 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33224 \$16 \$7545 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33226 \$153 \$9204 \$8614 \$9185 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33227 \$153 \$9293 \$9202 \$8898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33229 \$153 \$9139 \$9202 \$8728 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33230 \$153 \$9205 \$9202 \$8686 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33233 \$153 \$9205 \$8651 \$9185 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33234 \$16 \$8898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33235 \$16 \$8686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33236 \$16 \$8728 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33238 \$153 \$8899 \$9001 \$8890 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33239 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$33241 \$153 \$9162 \$9001 \$8647 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33244 \$153 \$9272 \$8818 \$8887 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33245 \$153 \$9162 \$8614 \$8887 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33246 \$16 \$9273 \$16 \$153 \$8635 VNB sky130_fd_sc_hd__clkbuf_2
X$33247 \$16 \$8647 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33248 \$153 \$9294 \$9001 \$8898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33249 \$153 \$9206 \$8277 \$9186 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33250 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$33252 \$16 \$8898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33253 \$153 \$9207 \$9001 \$8816 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33254 \$153 \$9207 \$8804 \$8887 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33255 \$153 \$9163 \$8651 \$8887 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33256 \$153 \$9274 \$8727 \$8887 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33257 \$16 \$8816 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33258 \$153 \$9164 \$9132 \$8686 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33261 \$153 \$9141 \$9132 \$8886 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33262 \$153 \$9208 \$8804 \$9111 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33263 \$16 \$8686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33264 \$153 \$9296 \$9132 \$8556 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33265 \$153 \$9164 \$8651 \$9111 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33267 \$153 \$9142 \$9132 \$8728 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33268 \$16 \$8556 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33269 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$33270 \$153 \$9247 \$9076 \$8886 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33271 \$153 \$9143 \$9076 \$8898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33273 \$153 \$9247 \$8727 \$9144 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33274 \$16 \$8898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33275 \$16 \$8728 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33276 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$33277 \$16 \$8886 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33278 \$16 \$7992 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33279 \$153 \$9225 \$9076 \$8556 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33281 \$153 \$9248 \$9076 \$8728 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33283 \$153 \$9225 \$8610 \$9144 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33284 \$153 \$9248 \$8818 \$9144 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33285 \$16 \$8556 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33286 \$16 \$6909 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33287 \$153 \$9297 \$9077 \$8886 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33288 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$33289 \$153 \$9145 \$9077 \$8898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33291 \$16 \$8886 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33293 \$153 \$9209 \$8804 \$9146 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33294 \$16 \$8898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33296 \$153 \$9249 \$9077 \$8890 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33297 \$153 \$9078 \$8610 \$9146 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33299 \$16 \$8890 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33300 \$153 \$9249 \$8277 \$9146 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33303 \$153 \$9165 \$8614 \$9146 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33305 \$153 \$9211 \$9044 \$8886 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33307 \$153 \$9226 \$9044 \$8890 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33308 \$16 \$8686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33309 \$16 \$8886 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33311 \$153 \$9210 \$8614 \$8989 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33312 \$16 \$8890 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33314 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$33315 \$153 \$9299 \$9044 \$8898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33316 \$153 \$9211 \$8727 \$8989 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33318 \$153 \$9212 \$8804 \$8989 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33319 \$16 \$8898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33320 \$16 \$8816 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33321 \$16 \$7072 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33323 \$16 \$8556 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33325 \$153 \$153 \$8727 \$9010 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33326 \$16 \$7288 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33327 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$33328 \$16 \$7065 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33329 \$153 \$153 \$8789 \$9010 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33330 \$153 \$153 \$8818 \$9010 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33331 \$153 \$153 \$8614 \$9010 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33332 \$153 \$9491 \$8818 \$9300 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33333 \$16 \$9227 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33334 \$16 \$7482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33335 \$153 \$9228 \$9116 \$9031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33337 \$153 \$8521 \$9116 \$9275 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33338 \$16 \$9031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33339 \$153 \$8751 \$9116 \$9253 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33340 \$16 \$9275 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33341 \$153 \$9213 \$8842 \$8126 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33343 \$16 \$7066 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33344 \$16 \$6582 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33345 \$153 \$9250 \$9116 \$9188 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33346 \$16 \$9253 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33347 \$153 \$9148 \$9116 \$9214 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33348 \$16 \$9188 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33349 \$16 \$8126 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33350 \$16 \$9214 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33351 \$16 \$7793 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33352 \$153 \$9187 \$9133 \$9324 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33353 \$16 \$9275 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33355 \$16 \$9045 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33356 \$16 \$9188 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33357 \$153 \$9251 \$8935 \$9275 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33358 \$153 \$9229 \$8935 \$9188 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33359 \$16 \$9031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33361 \$153 \$9251 \$9278 \$8958 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33362 \$16 \$8819 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33363 \$16 \$7484 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33366 \$153 \$9080 \$9047 \$8958 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33367 \$153 \$9261 \$9252 \$8958 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33369 \$16 \$7350 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33370 \$153 \$9168 \$9133 \$8958 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33371 \$16 \$9214 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33372 \$153 \$9169 \$8900 \$9214 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33373 \$16 \$9275 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33374 \$16 \$7903 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33375 \$16 \$7709 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33376 \$16 \$7668 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33378 \$16 \$7551 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33379 \$153 \$9169 \$9047 \$8891 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33380 \$16 \$7350 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33381 \$16 \$9253 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33382 \$153 \$9262 \$9252 \$8891 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33383 \$16 \$7350 \$16 \$153 \$8891 VNB sky130_fd_sc_hd__inv_1
X$33384 \$16 \$9253 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33385 \$16 \$9275 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33386 \$16 \$9214 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33388 \$153 \$9215 \$8972 \$9275 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33389 \$153 \$9171 \$9133 \$8840 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33391 \$16 \$8807 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33392 \$16 \$9031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33393 \$153 \$9215 \$9278 \$8840 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33394 \$153 \$9170 \$9047 \$8840 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33396 \$153 \$9277 \$9047 \$9276 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33397 \$153 \$9230 \$8972 \$9253 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33398 \$16 \$9455 \$16 \$153 \$8819 VNB sky130_fd_sc_hd__clkbuf_2
X$33401 \$153 \$9230 \$9252 \$8840 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33402 \$153 \$9172 \$8972 \$9188 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33404 \$153 \$9254 \$8937 \$9214 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33405 \$153 \$9172 \$8917 \$8840 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33409 \$153 \$9254 \$9047 \$8843 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33410 \$153 \$9189 \$8937 \$9188 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33411 \$16 \$9188 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33412 \$16 \$9188 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33413 \$153 \$9303 \$9050 \$9188 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33414 \$153 \$9083 \$9133 \$8843 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33415 \$153 \$9189 \$8917 \$8843 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33417 \$16 \$8869 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33418 \$16 \$7667 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33420 \$16 \$9275 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33421 \$16 \$8819 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33422 \$153 \$9255 \$9050 \$9275 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33423 \$16 \$7667 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33424 \$16 \$9045 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33425 \$153 \$9173 \$9050 \$9045 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33426 \$153 \$9255 \$9278 \$8993 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33428 \$153 \$9173 \$9174 \$8993 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33429 \$16 \$7952 \$8960 \$9305 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$33431 \$16 \$7540 \$8960 \$9149 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$33432 \$16 \$9214 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33433 \$153 \$9306 \$9052 \$9214 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33435 \$153 \$9032 \$9052 \$9031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33437 \$153 \$9216 \$9052 \$9253 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33438 \$16 \$9253 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33440 \$153 \$9084 \$9174 \$9033 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33441 \$16 \$7952 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33442 \$153 \$9326 \$9278 \$9033 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33443 \$153 \$9216 \$9252 \$9033 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33444 \$16 \$7540 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33445 \$16 \$7540 \$16 \$153 \$9033 VNB sky130_fd_sc_hd__inv_1
X$33447 \$16 \$7540 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33448 \$153 \$9118 \$8676 \$9033 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33449 \$16 \$9275 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33450 \$153 \$9307 \$9053 \$9275 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33451 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$33452 \$16 \$9031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33453 \$153 \$9176 \$9053 \$9031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33454 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$33455 \$16 \$9253 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33456 \$16 \$9188 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33458 \$153 \$9346 \$9053 \$9188 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33459 \$153 \$9176 \$9133 \$8920 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33460 \$153 \$9231 \$9054 \$9188 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33462 \$153 \$9217 \$9054 \$9253 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33464 \$16 \$9045 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33466 \$153 \$9217 \$9252 \$9151 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33467 \$153 \$9327 \$9347 \$9188 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33468 \$153 \$9347 \$7306 \$9232 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$33469 \$16 \$7431 \$8960 \$9232 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$33470 \$16 \$8936 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33471 \$153 \$9233 \$9054 \$9275 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33473 \$153 \$9309 \$9347 \$8936 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33474 \$153 \$9233 \$9278 \$9151 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33475 \$16 \$7431 \$16 \$153 \$9328 VNB sky130_fd_sc_hd__inv_1
X$33477 \$153 \$9234 \$9122 \$9152 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33478 \$16 \$9275 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33479 \$16 \$9055 \$8136 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$33481 \$16 \$7386 \$8824 \$9178 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$33482 \$153 \$9263 \$9059 \$9152 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33484 \$153 \$9234 \$9179 \$9134 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33485 \$153 \$9120 \$9179 \$8927 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33486 \$153 \$9190 \$8965 \$9152 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33487 \$16 \$8927 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33489 \$153 \$9310 \$9179 \$9035 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33490 \$153 \$9089 \$9122 \$8892 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33491 \$153 \$9153 \$9179 \$8879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33492 \$153 \$9311 \$9179 \$9154 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33494 \$16 \$8879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33496 \$153 \$9090 \$9059 \$8892 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33497 \$153 \$9190 \$9179 \$8844 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33498 \$16 \$9154 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33500 \$153 \$9235 \$8922 \$9134 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33501 \$16 \$8844 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33502 \$16 \$9134 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33503 \$16 \$7344 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33504 \$16 \$7350 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33507 \$16 \$9154 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33509 \$153 \$9020 \$9256 \$8906 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33510 \$153 \$9236 \$8922 \$9154 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33511 \$153 \$9279 \$7551 \$9237 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$33512 \$16 \$7350 \$8824 \$9237 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$33514 \$16 \$9035 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33515 \$153 \$9236 \$9103 \$8906 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33517 \$153 \$9125 \$8812 \$9035 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33518 \$16 \$7350 \$16 \$153 \$9264 VNB sky130_fd_sc_hd__inv_1
X$33519 \$153 \$9377 \$9122 \$9264 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33520 \$16 \$9191 \$16 \$153 \$8824 VNB sky130_fd_sc_hd__clkbuf_2
X$33521 \$153 \$9257 \$9256 \$9264 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33522 \$153 \$9123 \$8812 \$9134 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33524 \$153 \$9257 \$9279 \$8927 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33526 \$16 \$8893 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33528 \$153 \$9180 \$8874 \$9034 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33529 \$16 \$9034 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33530 \$16 \$8927 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33531 \$16 \$8383 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33533 \$153 \$9258 \$9279 \$8879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33536 \$153 \$9180 \$9059 \$8943 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33537 \$153 \$9155 \$8874 \$9134 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33539 \$153 \$9258 \$8923 \$9264 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33540 \$16 \$8879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33542 \$16 \$9034 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33543 \$153 \$9181 \$9103 \$8943 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33545 \$153 \$9315 \$8926 \$9034 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33547 \$16 \$8927 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33548 \$16 \$9154 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33549 \$153 \$8848 \$8926 \$8927 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33551 \$153 \$9058 \$8926 \$9154 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33553 \$153 \$9182 \$8977 \$8846 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33554 \$153 \$9281 \$9122 \$9280 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33556 \$16 \$9154 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33557 \$16 \$7540 \$8825 \$9238 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$33558 \$153 \$9316 \$7693 \$9238 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$33559 \$153 \$9093 \$8908 \$9154 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33561 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$33562 \$153 \$9094 \$8908 \$9134 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33564 \$153 \$9265 \$8977 \$9280 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33565 \$153 \$9259 \$9316 \$8844 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33566 \$16 \$7540 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33567 \$16 \$7540 \$16 \$153 \$9239 VNB sky130_fd_sc_hd__inv_1
X$33570 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$33571 \$153 \$9259 \$8965 \$9239 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33572 \$16 \$9134 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33573 \$153 \$8851 \$8877 \$9134 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33575 \$16 \$7306 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33576 \$153 \$9240 \$7306 \$9156 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$33577 \$153 \$9183 \$9103 \$8852 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33579 \$16 \$9034 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33580 \$153 \$9060 \$8877 \$9034 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33581 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$33582 \$16 \$8879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33583 \$153 \$9318 \$9240 \$8879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33585 \$153 \$9218 \$8996 \$9192 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33586 \$16 \$7431 \$16 \$153 \$9192 VNB sky130_fd_sc_hd__inv_1
X$33587 \$16 \$9134 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33589 \$153 \$9241 \$9240 \$8927 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33590 \$16 \$9134 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33591 \$153 \$9319 \$9240 \$9134 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33592 \$153 \$9241 \$9256 \$9192 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33593 \$153 \$9282 \$9059 \$9192 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33594 \$16 \$9035 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33595 \$153 \$9242 \$9240 \$9035 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33598 \$153 \$9320 \$9240 \$9154 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33599 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$33600 \$153 \$9242 \$8977 \$9192 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33601 \$153 \$9184 \$9059 \$8947 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33602 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$33604 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$33605 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$33606 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$33607 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$33608 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$33609 \$153 \$5175 \$5174 \$4579 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33611 \$16 \$4579 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33612 \$153 \$5225 \$5266 \$5181 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33613 \$153 \$5225 \$5174 \$5120 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33614 \$153 \$5021 \$4864 \$3385 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33615 \$16 \$5181 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33616 \$16 \$3616 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33618 \$16 \$3692 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33621 \$16 \$5736 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33622 \$16 \$3385 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33623 \$153 \$5313 \$5266 \$5274 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33624 \$153 \$4864 \$5226 \$5121 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$33625 \$16 \$5274 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33627 \$16 \$3692 \$5176 \$5164 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$33629 \$153 \$4968 \$3307 \$4859 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33631 \$153 \$5266 \$5151 \$5164 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$33633 \$153 \$5239 \$5200 \$5181 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33635 \$153 \$5165 \$5177 \$4579 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33636 \$16 \$5226 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33637 \$16 \$5176 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33638 \$153 \$5178 \$5463 \$5166 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33639 \$16 \$4893 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33641 \$153 \$5239 \$5174 \$5166 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33642 \$153 \$5200 \$3767 \$5179 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$33643 \$153 \$5315 \$5200 \$5245 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33644 \$153 \$5180 \$5055 \$5166 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33645 \$16 \$3841 \$5176 \$5179 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$33647 \$153 \$5148 \$4614 \$3571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33648 \$16 \$5245 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33650 \$153 \$5227 \$5240 \$5274 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33651 \$153 \$5148 \$3422 \$4707 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33652 \$16 \$3571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33653 \$16 \$3778 \$5176 \$5241 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$33654 \$153 \$5149 \$4789 \$3571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33656 \$153 \$5240 \$4079 \$5241 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$33657 \$153 \$5149 \$3422 \$4693 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33658 \$153 \$5275 \$5055 \$5276 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33660 \$16 \$4896 \$4538 \$5023 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$33662 \$153 \$5242 \$5267 \$5274 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33664 \$153 \$5105 \$3389 \$4693 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33665 \$16 \$4538 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33666 \$16 \$4896 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33667 \$153 \$5242 \$4706 \$5277 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33668 \$153 \$5167 \$4865 \$3385 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33670 \$16 \$3714 \$5176 \$5278 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$33673 \$153 \$5167 \$3394 \$4940 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33674 \$153 \$5243 \$5267 \$5181 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33675 \$16 \$3385 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33676 \$153 \$4865 \$4973 \$5122 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$33677 \$153 \$5243 \$5174 \$5277 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33679 \$16 \$5181 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33680 \$153 \$5244 \$5347 \$5181 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33682 \$153 \$5123 \$3389 \$4940 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33684 \$153 \$5182 \$5107 \$5168 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33685 \$153 \$5244 \$5174 \$5168 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33687 \$153 \$5054 \$5347 \$5736 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33688 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$33691 \$16 \$3761 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33692 \$16 \$3761 \$16 \$153 \$5168 VNB sky130_fd_sc_hd__inv_1
X$33693 \$153 \$5279 \$4706 \$5168 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33694 \$16 \$5736 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33696 \$153 \$4867 \$5109 \$5124 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$33698 \$153 \$5316 \$5246 \$5245 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33699 \$16 \$3616 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33701 \$16 \$5109 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33703 \$16 \$5245 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33705 \$16 \$5181 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33706 \$153 \$5150 \$4791 \$3571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33707 \$153 \$5280 \$5246 \$5181 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33708 \$153 \$5150 \$3422 \$4941 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33710 \$16 \$3997 \$16 \$153 \$5337 VNB sky130_fd_sc_hd__inv_1
X$33711 \$16 \$3997 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33714 \$16 \$5184 \$3660 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$33715 \$153 \$5053 \$3394 \$4359 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33716 \$16 \$5184 \$3767 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$33717 \$16 \$5268 \$5226 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$33718 \$16 \$5268 \$5314 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$33719 \$16 \$5184 \$5183 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$33720 \$16 \$5268 \$4973 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$33721 \$16 \$5268 \$4939 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$33722 \$16 \$5184 \$4079 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$33723 \$16 \$5281 \$16 \$153 \$5268 VNB sky130_fd_sc_hd__clkbuf_2
X$33724 \$16 \$5184 \$5151 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$33725 \$16 \$5281 \$16 \$153 \$5184 VNB sky130_fd_sc_hd__clkbuf_2
X$33726 \$16 \$5184 \$4083 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$33727 \$16 \$3907 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33728 \$16 \$4869 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33729 \$16 \$5269 \$4616 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$33731 \$16 \$5184 \$5201 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$33732 \$16 \$5281 \$16 \$153 \$5269 VNB sky130_fd_sc_hd__clkbuf_2
X$33733 \$16 \$5106 \$3949 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$33734 \$16 \$3906 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33735 \$153 \$4711 \$4943 \$5202 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$33736 \$16 \$4822 \$4012 \$5202 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$33737 \$16 \$1482 \$16 \$153 \$5281 VNB sky130_fd_sc_hd__clkbuf_2
X$33738 \$16 \$5281 \$16 \$153 \$5106 VNB sky130_fd_sc_hd__clkbuf_2
X$33739 \$16 \$5106 \$3906 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$33740 \$16 \$5106 \$4246 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$33741 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33742 \$16 \$5106 \$5228 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$33743 \$153 \$5126 \$3389 \$4694 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33744 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33746 \$153 \$153 \$5174 \$5203 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33748 \$16 \$4620 \$16 \$153 \$5203 VNB sky130_fd_sc_hd__clkbuf_2
X$33749 \$153 \$3865 \$1482 \$4706 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33751 \$153 \$3633 \$1482 \$5177 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33752 \$16 \$5177 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33754 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33755 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33757 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33759 \$153 \$3952 \$1482 \$5174 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33760 \$153 \$3617 \$1482 \$5055 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33761 \$16 \$5174 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33762 \$16 \$3778 \$5186 \$5127 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$33764 \$16 \$4978 \$16 \$153 \$4896 VNB sky130_fd_sc_hd__clkbuf_2
X$33765 \$16 \$5055 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33766 \$16 \$5226 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33768 \$16 \$4902 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33771 \$16 \$5152 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33772 \$153 \$5185 \$5128 \$5271 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33773 \$153 \$4926 \$5152 \$5060 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$33774 \$153 \$5185 \$5069 \$5169 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33775 \$16 \$3778 \$16 \$153 \$5169 VNB sky130_fd_sc_hd__inv_1
X$33776 \$16 \$5271 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33778 \$153 \$5187 \$5128 \$5232 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33781 \$16 \$5186 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33782 \$16 \$5186 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33783 \$16 \$3692 \$5186 \$5204 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$33784 \$153 \$5187 \$5205 \$5169 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33785 \$153 \$5248 \$5151 \$5204 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$33787 \$153 \$5029 \$4926 \$3480 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33788 \$16 \$3778 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33791 \$153 \$5249 \$5248 \$5232 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33792 \$16 \$3480 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33793 \$16 \$5080 \$4275 \$5188 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$33794 \$153 \$4873 \$5051 \$5188 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$33795 \$16 \$3692 \$16 \$153 \$5270 VNB sky130_fd_sc_hd__inv_1
X$33796 \$153 \$5250 \$5248 \$5271 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33799 \$153 \$5108 \$4873 \$3543 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33800 \$153 \$5251 \$5248 \$5324 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33801 \$16 \$3543 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33802 \$153 \$5034 \$4873 \$3480 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33803 \$16 \$4896 \$4275 \$5229 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$33805 \$153 \$5350 \$3767 \$5282 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$33806 \$153 \$5189 \$5205 \$5013 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33807 \$16 \$4275 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33808 \$153 \$5206 \$5096 \$5013 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33809 \$16 \$5095 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33810 \$153 \$5253 \$5095 \$5252 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$33812 \$16 \$3761 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33814 \$16 \$3761 \$5186 \$5252 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$33815 \$16 \$4893 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33816 \$16 \$5314 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33817 \$16 \$5186 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33818 \$153 \$4622 \$5314 \$5129 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$33819 \$153 \$5319 \$5253 \$5271 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33820 \$153 \$5061 \$3354 \$4818 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33821 \$16 \$3761 \$16 \$153 \$5170 VNB sky130_fd_sc_hd__inv_1
X$33824 \$16 \$3543 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33825 \$153 \$5190 \$5096 \$5170 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33826 \$153 \$5320 \$5253 \$5232 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33828 \$16 \$4973 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33829 \$153 \$4875 \$4973 \$5130 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$33830 \$16 \$3714 \$5186 \$5272 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$33831 \$16 \$5232 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33832 \$153 \$5321 \$5231 \$5232 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33834 \$153 \$5191 \$5209 \$5170 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33835 \$16 \$3714 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33836 \$16 \$5338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33837 \$153 \$5207 \$5231 \$5338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33838 \$16 \$3714 \$16 \$153 \$5283 VNB sky130_fd_sc_hd__inv_1
X$33839 \$16 \$5232 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33841 \$153 \$5284 \$5096 \$5283 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33843 \$153 \$5153 \$4875 \$3480 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33844 \$153 \$5322 \$5069 \$5283 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33846 \$153 \$5285 \$5254 \$5232 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33847 \$153 \$5153 \$3504 \$4798 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33848 \$16 \$3480 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33849 \$16 \$5232 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33851 \$16 \$5109 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33852 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$33853 \$153 \$5037 \$4876 \$3480 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33854 \$153 \$5255 \$5254 \$5271 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33855 \$153 \$5208 \$5209 \$5171 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33856 \$153 \$5255 \$5069 \$5171 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33857 \$153 \$5131 \$3556 \$4696 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33859 \$16 \$3480 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33861 \$153 \$5256 \$5273 \$5232 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33862 \$16 \$3543 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33864 \$153 \$4948 \$4943 \$5132 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$33865 \$153 \$5256 \$5205 \$5286 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33866 \$16 \$3886 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33869 \$153 \$5154 \$4948 \$3543 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33870 \$153 \$5257 \$5273 \$5271 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33871 \$153 \$5257 \$5069 \$5286 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33872 \$153 \$5154 \$3556 \$5066 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33873 \$16 \$3543 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33875 \$16 \$16 \$153 VNB sky130_fd_sc_hd__conb_1
X$33878 \$16 \$5271 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33879 \$16 \$4620 \$16 \$153 \$5155 VNB sky130_fd_sc_hd__clkbuf_2
X$33880 \$16 \$3344 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33881 \$153 \$153 \$5069 \$5155 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33882 \$153 \$153 \$5287 \$5155 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33883 \$153 \$153 \$5390 \$5155 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33884 \$153 \$153 \$5205 \$5155 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33885 \$153 \$153 \$5406 \$5155 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33886 \$16 \$4620 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33888 \$16 \$5390 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33890 \$16 \$5205 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33891 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33894 \$153 \$4049 \$1482 \$5519 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33895 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33896 \$153 \$3598 \$1482 \$5390 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33897 \$16 \$5324 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33898 \$16 \$5287 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33899 \$153 \$4984 \$3435 \$5066 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33900 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33901 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33903 \$153 \$4408 \$1482 \$5287 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33904 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$33905 \$16 \$3889 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33906 \$153 \$5211 \$5110 \$3889 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33908 \$153 \$5288 \$5110 \$3960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33910 \$153 \$5133 \$3858 \$4801 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33911 \$153 \$5233 \$5110 \$3792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33913 \$153 \$5233 \$3939 \$5172 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33914 \$153 \$5212 \$5110 \$3791 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33915 \$16 \$3792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33916 \$16 \$4760 \$4881 \$5289 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$33918 \$153 \$5326 \$5110 \$3814 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33919 \$153 \$5134 \$3763 \$5172 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33921 \$16 \$3791 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33923 \$16 \$3792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33924 \$153 \$5070 \$3788 \$5015 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33925 \$153 \$5111 \$5039 \$3792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33927 \$153 \$5213 \$5039 \$3791 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33928 \$16 \$3814 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33929 \$16 \$4930 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33930 \$16 \$4834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33931 \$153 \$5290 \$3716 \$5015 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33932 \$153 \$5213 \$3919 \$5015 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33933 \$16 \$4834 \$16 \$153 \$5015 VNB sky130_fd_sc_hd__inv_1
X$33934 \$16 \$3791 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33936 \$16 \$3792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33937 \$153 \$5156 \$5041 \$3791 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33939 \$153 \$5258 \$5041 \$3792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33941 \$153 \$5156 \$3919 \$5016 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33942 \$153 \$5258 \$3939 \$5016 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33943 \$16 \$3792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33946 \$153 \$5234 \$5042 \$3792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33948 \$153 \$5214 \$5042 \$3814 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33949 \$153 \$5291 \$3651 \$5016 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33950 \$153 \$5234 \$3939 \$4951 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33951 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$33952 \$16 \$4949 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33953 \$16 \$4048 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33954 \$16 \$3731 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33956 \$153 \$5292 \$5042 \$4048 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33957 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$33959 \$16 \$5331 \$16 \$153 \$4951 VNB sky130_fd_sc_hd__inv_1
X$33960 \$16 \$5331 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33962 \$153 \$5192 \$3716 \$4951 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33964 \$16 \$5498 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33965 \$16 \$3792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33966 \$16 \$5017 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33967 \$153 \$5260 \$4931 \$3792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33968 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$33971 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$33972 \$16 \$3814 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33973 \$153 \$5136 \$3919 \$4992 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33974 \$153 \$5260 \$3939 \$4992 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33975 \$16 \$3791 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33976 \$153 \$5293 \$3651 \$4992 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33977 \$16 \$3852 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33978 \$153 \$5215 \$4952 \$3814 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33981 \$153 \$5294 \$4952 \$3792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33982 \$16 \$3792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33983 \$16 \$4724 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33984 \$153 \$5137 \$3919 \$5138 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33985 \$153 \$5294 \$3939 \$5138 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33986 \$16 \$4882 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33987 \$16 \$4882 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33988 \$16 \$3792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33989 \$16 \$3791 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33991 \$153 \$5295 \$4920 \$3792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$33992 \$153 \$4993 \$3788 \$5138 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33993 \$16 \$5353 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33994 \$16 \$5216 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33995 \$16 \$5158 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33996 \$16 \$4885 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$33997 \$153 \$5295 \$3939 \$4953 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33998 \$153 \$5193 \$3651 \$4953 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$33999 \$16 \$5354 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34000 \$16 \$3792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34002 \$16 \$4954 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34004 \$16 \$5400 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34005 \$153 \$5261 \$5043 \$3792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34006 \$16 \$5173 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34007 \$16 \$5173 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34008 \$153 \$4996 \$3788 \$5139 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34009 \$153 \$5090 \$3919 \$5139 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34010 \$153 \$5261 \$3939 \$5139 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34011 \$16 \$3960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34014 \$153 \$5296 \$5112 \$3960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34016 \$153 \$5217 \$5112 \$3792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34017 \$153 \$5112 \$5235 \$5262 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$34018 \$16 \$5173 \$16 \$153 \$5113 VNB sky130_fd_sc_hd__inv_1
X$34019 \$153 \$5218 \$5112 \$3731 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34021 \$16 \$5173 \$4724 \$5262 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$34022 \$153 \$5263 \$5112 \$4048 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34023 \$153 \$5218 \$3788 \$5113 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34024 \$16 \$5194 \$4609 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$34025 \$153 \$4543 \$4414 \$5158 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34026 \$153 \$5263 \$3858 \$5113 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34028 \$153 \$4885 \$3719 \$4954 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34030 \$153 \$5216 \$3565 \$5158 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34031 \$153 \$5157 \$4912 \$4935 \$4933 \$4833 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$34032 \$153 \$4933 \$4833 \$5297 \$4912 \$4935 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$34033 \$153 \$4912 \$4933 \$5219 \$4833 \$4935 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$34034 \$16 \$5219 \$16 \$153 \$5259 VNB sky130_fd_sc_hd__clkbuf_2
X$34035 \$16 \$5355 \$5264 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$34036 \$16 \$5157 \$16 \$153 \$4760 VNB sky130_fd_sc_hd__clkbuf_2
X$34038 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34039 \$16 \$4834 \$5116 \$5298 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$34041 \$153 \$5195 \$5001 \$4936 \$4937 \$4958 \$16 \$16 VNB
+ sky130_fd_sc_hd__nor4b_2
X$34042 \$153 \$4936 \$4937 \$5300 \$5001 \$4958 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$34043 \$153 \$5196 \$5452 \$5299 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$34044 \$153 \$5001 \$4937 \$5220 \$4936 \$4958 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$34045 \$16 \$5806 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34047 \$153 \$5159 \$5196 \$3721 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34048 \$16 \$3826 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34049 \$153 \$5142 \$5196 \$4057 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34050 \$153 \$5159 \$3676 \$5114 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34051 \$16 \$5220 \$16 \$153 \$5173 VNB sky130_fd_sc_hd__clkbuf_2
X$34052 \$16 \$5300 \$16 \$153 \$5400 VNB sky130_fd_sc_hd__clkbuf_2
X$34054 \$153 \$5160 \$5196 \$3680 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34056 \$153 \$5115 \$5196 \$3602 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34057 \$153 \$5160 \$3719 \$5114 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34058 \$153 \$5301 \$3142 \$5114 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34059 \$16 \$4760 \$16 \$153 \$5114 VNB sky130_fd_sc_hd__inv_1
X$34061 \$16 \$3680 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34062 \$16 \$3826 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34064 \$16 \$3680 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34065 \$153 \$4961 \$5197 \$4057 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34067 \$153 \$5302 \$3986 \$5019 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34068 \$153 \$5100 \$5197 \$3602 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34070 \$153 \$5161 \$5197 \$3721 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34072 \$16 \$3602 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34073 \$153 \$5161 \$3676 \$5019 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34074 \$16 \$3721 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34075 \$16 \$4057 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34077 \$16 \$3680 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34078 \$16 \$3691 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34079 \$153 \$5101 \$5303 \$3680 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34080 \$16 \$5259 \$16 \$153 \$5117 VNB sky130_fd_sc_hd__inv_1
X$34081 \$153 \$5143 \$5303 \$3602 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34083 \$16 \$5259 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34084 \$16 \$5017 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34085 \$16 \$3602 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34086 \$16 \$3567 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34087 \$16 \$3721 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34088 \$16 \$4057 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34089 \$153 \$5221 \$5303 \$3721 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34090 \$153 \$5118 \$5303 \$4057 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34091 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$34093 \$16 \$4057 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34095 \$16 \$3721 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34096 \$153 \$5102 \$5198 \$4057 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34097 \$153 \$5162 \$5198 \$3721 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34098 \$153 \$5304 \$3986 \$5119 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34099 \$153 \$5162 \$3676 \$5119 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34102 \$153 \$5265 \$3676 \$3567 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34104 \$153 \$5222 \$5198 \$3602 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34105 \$153 \$5222 \$3565 \$5119 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34106 \$153 \$4997 \$5163 \$3721 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34107 \$153 \$5305 \$3860 \$5119 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34108 \$16 \$5400 \$16 \$153 \$4954 VNB sky130_fd_sc_hd__inv_1
X$34110 \$153 \$4916 \$3860 \$5011 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34111 \$153 \$5223 \$5163 \$3602 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34112 \$153 \$4782 \$5163 \$4057 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34113 \$16 \$3680 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34114 \$16 \$3602 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34115 \$16 \$4057 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34116 \$153 \$4764 \$3142 \$5011 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34117 \$16 \$5473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34119 \$16 \$5173 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34120 \$16 \$5235 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34121 \$16 \$3721 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34122 \$153 \$4461 \$5144 \$3721 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34123 \$153 \$4543 \$5144 \$4057 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34125 \$16 \$4057 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34126 \$16 \$3602 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34127 \$16 \$5354 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34128 \$153 \$5216 \$5144 \$3602 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34129 \$16 \$5306 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34132 \$16 \$5002 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34133 \$16 \$5173 \$4736 \$5237 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$34134 \$153 \$5224 \$4414 \$4965 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34135 \$153 \$4892 \$5235 \$5237 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$34136 \$153 \$5307 \$3142 \$4965 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34137 \$153 \$5308 \$4892 \$3691 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34140 \$153 \$5103 \$5199 \$3680 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34141 \$16 \$5173 \$16 \$153 \$4963 VNB sky130_fd_sc_hd__inv_1
X$34142 \$153 \$4966 \$5199 \$3602 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34143 \$16 \$3602 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34144 \$153 \$5310 \$5074 \$5309 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34146 \$16 \$5354 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34147 \$16 \$3721 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34149 \$153 \$5046 \$5199 \$3721 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34150 \$153 \$5224 \$5199 \$4057 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34151 \$16 \$5173 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34152 \$16 \$4057 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34153 \$153 \$5311 \$5509 \$5309 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34154 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$34157 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$34158 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$34159 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$34160 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$34161 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$34162 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$34163 \$153 \$10135 \$10427 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$34164 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$34166 \$153 \$10398 \$10256 \$10427 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34167 \$16 \$10135 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34169 \$16 \$10427 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34170 \$153 \$10398 \$10327 \$10245 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34173 \$153 \$10329 \$10256 \$10646 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34174 \$153 \$10410 \$10256 \$10367 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34175 \$16 \$10646 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34177 \$153 \$10410 \$10330 \$10245 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34178 \$16 \$10367 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34179 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$34181 \$153 \$10411 \$10256 \$10476 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34182 \$16 \$10348 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34183 \$16 \$10348 \$16 \$153 \$10245 VNB sky130_fd_sc_hd__inv_1
X$34184 \$153 \$10256 \$10603 \$10488 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$34186 \$153 \$10347 \$10250 \$10295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34187 \$16 \$10348 \$10468 \$10488 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$34189 \$16 \$10427 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34191 \$153 \$10428 \$10250 \$10427 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34192 \$16 \$10476 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34193 \$16 \$10295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34194 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$34195 \$153 \$10257 \$10250 \$10646 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34196 \$153 \$10377 \$10250 \$10476 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34198 \$153 \$10377 \$10705 \$10210 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34199 \$16 \$10539 \$16 \$153 \$10210 VNB sky130_fd_sc_hd__inv_1
X$34200 \$16 \$10476 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34203 \$153 \$10258 \$10251 \$10646 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34204 \$153 \$10399 \$10251 \$10367 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34205 \$153 \$10399 \$10330 \$10211 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34206 \$16 \$10367 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34209 \$16 \$10453 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34210 \$16 \$10453 \$10468 \$10469 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$34211 \$16 \$10646 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34213 \$153 \$10429 \$10251 \$10476 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34214 \$16 \$10427 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34215 \$153 \$10454 \$10251 \$10427 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34216 \$153 \$10454 \$10327 \$10211 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34218 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$34219 \$16 \$10476 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34220 \$16 \$10427 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34221 \$153 \$10430 \$10259 \$10646 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34222 \$153 \$10412 \$10259 \$10427 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34223 \$16 \$10646 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34224 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$34225 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$34227 \$153 \$10350 \$10259 \$10295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34228 \$153 \$10412 \$10327 \$10246 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34229 \$153 \$10430 \$10318 \$10246 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34230 \$153 \$10350 \$10276 \$10246 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34232 \$153 \$10378 \$10199 \$10427 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34233 \$16 \$10295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34236 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$34237 \$153 \$10378 \$10327 \$10212 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34238 \$153 \$10490 \$10199 \$10646 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34239 \$16 \$6693 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34240 \$16 \$10368 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34241 \$16 \$10226 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34242 \$16 \$10413 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34243 \$153 \$8838 \$10367 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$34244 \$16 \$10367 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34245 \$16 \$10646 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34248 \$16 \$10295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34250 \$16 \$10295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34251 \$153 \$10143 \$10476 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$34252 \$153 \$9898 \$8209 \$9866 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34253 \$16 \$8838 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34254 \$16 \$10143 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34255 \$153 \$10431 \$10252 \$10476 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34257 \$153 \$10455 \$10252 \$10427 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34258 \$153 \$10455 \$10327 \$10331 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34259 \$153 \$10332 \$10252 \$10368 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34260 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$34263 \$153 \$10432 \$10456 \$10226 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34264 \$153 \$10333 \$10252 \$10646 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34265 \$153 \$9227 \$10646 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$34266 \$16 \$9227 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34267 \$16 \$10368 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34268 \$16 \$10646 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34271 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$34273 \$16 \$8638 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34274 \$153 \$10351 \$10456 \$10295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34275 \$16 \$10318 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34276 \$16 \$10330 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34277 \$153 \$9869 \$10295 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$34279 \$16 \$9869 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34281 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34282 \$153 \$10144 \$8340 \$10705 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34283 \$153 \$10201 \$8340 \$10330 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34284 \$153 \$10433 \$8340 \$10327 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34285 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34286 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34288 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34290 \$153 \$10146 \$8340 \$10161 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34291 \$16 \$10327 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34293 \$153 \$10379 \$10320 \$10606 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34294 \$16 \$10260 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34295 \$16 \$10348 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34296 \$153 \$10379 \$10344 \$10369 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34297 \$16 \$10348 \$16 \$153 \$10369 VNB sky130_fd_sc_hd__inv_1
X$34299 \$153 \$10457 \$10516 \$10369 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34300 \$153 \$10352 \$10320 \$10338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34301 \$153 \$10458 \$10686 \$10369 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34302 \$153 \$10352 \$10309 \$10369 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34303 \$16 \$10319 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34304 \$153 \$10494 \$10320 \$10470 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34305 \$16 \$10338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34307 \$153 \$10335 \$10320 \$10382 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34308 \$153 \$10353 \$10401 \$10369 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34309 \$16 \$10298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34310 \$153 \$10459 \$10247 \$10477 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34311 \$153 \$10460 \$10400 \$10338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34312 \$16 \$10470 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34315 \$153 \$10460 \$10309 \$10337 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34316 \$16 \$10338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34317 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$34319 \$153 \$10354 \$10400 \$10298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34320 \$153 \$10434 \$10400 \$10606 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34322 \$153 \$10434 \$10344 \$10337 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34323 \$153 \$10354 \$10401 \$10337 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34324 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$34325 \$16 \$10606 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34327 \$153 \$10495 \$10380 \$10606 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34328 \$153 \$10355 \$10380 \$10338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34330 \$153 \$10496 \$10380 \$10470 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34331 \$16 \$10338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34332 \$16 \$10606 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34333 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$34334 \$153 \$10414 \$10380 \$10382 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34335 \$16 \$10470 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34336 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$34337 \$153 \$10414 \$10098 \$10339 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34338 \$16 \$10382 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34340 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$34342 \$153 \$10498 \$10381 \$10606 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34343 \$153 \$10356 \$10381 \$10338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34344 \$16 \$10606 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34346 \$16 \$10555 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34347 \$153 \$10402 \$10381 \$10298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34348 \$16 \$8890 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34351 \$153 \$10435 \$10381 \$10382 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34352 \$153 \$10402 \$10401 \$10515 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34353 \$16 \$10382 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34354 \$16 \$10470 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34355 \$16 \$10298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34357 \$16 \$8607 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34358 \$16 \$10322 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34359 \$153 \$10248 \$10340 \$10470 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34360 \$16 \$8411 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34362 \$153 \$10461 \$10340 \$10338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34363 \$153 \$10461 \$10309 \$10249 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34365 \$153 \$10415 \$10340 \$10298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34366 \$16 \$10338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34367 \$16 \$10470 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34368 \$16 \$10253 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34370 \$16 \$8555 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34371 \$153 \$10415 \$10401 \$10249 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34372 \$153 \$10341 \$10340 \$10382 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34373 \$16 \$10298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34374 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$34375 \$153 \$10436 \$10323 \$10514 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34376 \$16 \$10382 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34378 \$16 \$10262 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34379 \$16 \$10338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34382 \$153 \$10416 \$10323 \$10382 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34383 \$153 \$10436 \$10538 \$10343 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34384 \$153 \$10416 \$10098 \$10343 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34385 \$153 \$10358 \$10401 \$10343 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34386 \$16 \$10298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34387 \$16 \$10382 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34388 \$153 \$10403 \$10247 \$10343 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34391 \$153 \$10139 \$10514 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$34392 \$153 \$10068 \$8804 \$9845 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34393 \$153 \$9925 \$8614 \$9845 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34394 \$153 \$10238 \$10470 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$34396 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34398 \$153 \$10043 \$10338 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$34399 \$153 \$7949 \$7934 \$10500 \$7829 \$16 \$16 VNB
+ sky130_fd_sc_hd__nor3b_4
X$34400 \$153 \$9969 \$8610 \$9845 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34403 \$16 \$7949 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34405 \$153 \$9227 \$10300 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$34406 \$16 \$7949 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34407 \$16 \$7934 \$7949 \$7829 \$153 \$16 \$10478 VNB sky130_fd_sc_hd__and3_4
X$34408 \$153 \$10345 \$8340 \$10686 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34409 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34410 \$16 \$10043 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34411 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34413 \$153 \$8838 \$10578 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$34414 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34415 \$16 \$8838 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34417 \$16 \$10135 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34418 \$153 \$10135 \$10551 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$34419 \$153 \$8839 \$10386 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$34421 \$153 \$10260 \$8340 \$10471 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34422 \$153 \$10202 \$8340 \$10370 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34423 \$153 \$10147 \$8340 \$10472 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34425 \$153 \$10384 \$8340 \$10516 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34426 \$153 \$153 \$10501 \$10479 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34427 \$153 \$10462 \$10833 \$10480 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34429 \$153 \$6911 \$8347 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$34430 \$16 \$10578 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34431 \$16 \$10471 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34432 \$16 \$10417 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34434 \$16 \$10472 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34436 \$16 \$10386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34437 \$153 \$10371 \$10463 \$10386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34438 \$153 \$10280 \$9047 \$9871 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34439 \$153 \$10231 \$8917 \$9871 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34440 \$153 \$10464 \$10370 \$10372 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34443 \$153 \$10281 \$9252 \$9871 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34445 \$16 \$10386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34446 \$16 \$10300 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34447 \$153 \$10437 \$10528 \$10386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34448 \$16 \$6993 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34449 \$153 \$10360 \$8917 \$9953 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34450 \$153 \$6993 \$10311 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$34451 \$16 \$10473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34454 \$153 \$10481 \$10417 \$10482 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34455 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$34456 \$153 \$10371 \$10472 \$10372 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34457 \$16 \$10300 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34458 \$153 \$10385 \$10474 \$10300 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34459 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$34460 \$16 \$9253 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34464 \$153 \$10385 \$10417 \$10373 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34465 \$153 \$10465 \$10501 \$10372 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34466 \$16 \$6984 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34467 \$153 \$10483 \$10472 \$10373 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34468 \$153 \$6984 \$10361 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$34469 \$16 \$10473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34471 \$16 \$10473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34472 \$16 \$10578 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34475 \$153 \$10438 \$10404 \$10578 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34476 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$34477 \$16 \$10386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34478 \$153 \$10405 \$10404 \$10386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34479 \$153 \$10314 \$8917 \$10009 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34481 \$153 \$9776 \$9133 \$9642 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34483 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$34484 \$16 \$10300 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34485 \$16 \$10578 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34486 \$153 \$10406 \$10387 \$10578 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34488 \$153 \$10439 \$10387 \$10300 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34489 \$16 \$10386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34490 \$16 \$9642 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34491 \$153 \$10407 \$10387 \$10386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34492 \$16 \$10473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34494 \$153 \$10440 \$10387 \$10473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34495 \$153 \$10439 \$10417 \$10374 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34496 \$16 \$9642 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34497 \$16 \$10473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34498 \$16 \$10300 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34499 \$16 \$12245 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34500 \$153 \$10441 \$10475 \$10300 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34501 \$16 \$10597 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34504 \$16 \$10386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34506 \$16 \$9188 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34507 \$153 \$10389 \$10157 \$9188 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34508 \$153 \$10442 \$10475 \$10473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34509 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$34510 \$16 \$10473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34511 \$16 \$10386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34512 \$153 \$10362 \$10388 \$10473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34515 \$153 \$10443 \$10388 \$10386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34516 \$153 \$10389 \$8917 \$9872 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34517 \$16 \$10611 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34519 \$16 \$7115 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34521 \$153 \$7115 \$10383 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$34522 \$16 \$10277 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34524 \$153 \$10362 \$10501 \$10375 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34525 \$16 \$10345 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34526 \$153 \$10075 \$4303 \$10277 \$10345 \$10390 \$10391 \$10220 \$16 \$16
+ VNB sky130_fd_sc_hd__mux4_1
X$34528 \$16 \$9275 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34530 \$153 \$10315 \$10417 \$10375 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34532 \$16 \$10278 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34533 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34534 \$16 \$10384 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34535 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34536 \$16 \$10265 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34537 \$153 \$10266 \$8340 \$10560 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34538 \$16 \$10529 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34539 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34540 \$153 \$10159 \$8340 \$10376 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34541 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34542 \$153 \$10084 \$8340 \$10694 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34545 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34546 \$153 \$10204 \$8340 \$10285 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34547 \$153 \$10391 \$8340 \$9122 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34548 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34550 \$153 \$10527 \$10392 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$34552 \$16 \$9122 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34553 \$16 \$10408 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34554 \$153 \$10485 \$10466 \$10484 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34555 \$16 \$10238 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34556 \$153 \$10238 \$10326 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$34558 \$153 \$10286 \$9122 \$9981 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34559 \$16 \$10527 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34561 \$16 \$9256 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34562 \$16 \$10408 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34563 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$34564 \$153 \$7178 \$10527 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$34566 \$153 \$7095 \$10139 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$34567 \$16 \$7178 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34570 \$16 \$7095 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34571 \$16 \$10446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34572 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$34573 \$153 \$10205 \$10467 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$34575 \$153 \$7034 \$10043 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$34576 \$16 \$10205 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34577 \$16 \$11016 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34580 \$16 \$7034 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34581 \$153 \$10043 \$10393 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$34583 \$153 \$7098 \$9997 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$34584 \$153 \$9997 \$10446 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$34585 \$16 \$7098 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34586 \$16 \$9997 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34589 \$16 \$10393 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34590 \$153 \$10507 \$10444 \$10393 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34591 \$153 \$10288 \$9059 \$10011 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34592 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$34593 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$34594 \$153 \$10445 \$10444 \$10346 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34596 \$16 \$10097 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34598 \$153 \$10240 \$8923 \$10011 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34599 \$153 \$10289 \$9122 \$10011 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34600 \$153 \$10445 \$10285 \$10519 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34602 \$153 \$10487 \$10376 \$10519 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34603 \$16 \$10326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34604 \$16 \$10346 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34605 \$153 \$10418 \$10394 \$10346 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34607 \$153 \$10509 \$10394 \$10446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34608 \$153 \$10419 \$10394 \$10326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34609 \$153 \$10418 \$10285 \$10520 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34610 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$34613 \$16 \$10446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34614 \$16 \$10346 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34615 \$153 \$10447 \$10395 \$10446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34616 \$153 \$10420 \$10395 \$10346 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34617 \$153 \$10290 \$9059 \$9988 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34619 \$153 \$9917 \$9059 \$10222 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34620 \$153 \$9862 \$8977 \$10222 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34622 \$16 \$10222 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34623 \$16 \$10446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34624 \$16 \$10393 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34625 \$16 \$10346 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34626 \$153 \$10421 \$10325 \$10346 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34627 \$153 \$10448 \$10325 \$10446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34628 \$16 \$10222 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34631 \$16 \$10326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34634 \$16 \$10446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34635 \$16 \$10409 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34636 \$153 \$8479 \$7376 \$8429 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34637 \$16 \$10393 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34638 \$16 \$8429 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34639 \$153 \$10422 \$10396 \$10393 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34640 \$153 \$10450 \$10396 \$10326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34641 \$153 \$8085 \$7462 \$7076 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34644 \$16 \$10510 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34646 \$153 \$10449 \$10396 \$10446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34647 \$153 \$10423 \$10396 \$10346 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34648 \$16 \$10564 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34649 \$16 \$9034 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34651 \$16 \$7076 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34652 \$153 \$10114 \$8996 \$10112 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34654 \$16 \$10346 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34656 \$16 \$8055 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34657 \$153 \$10424 \$10397 \$10346 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34658 \$153 \$10451 \$10397 \$10326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34659 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$34660 \$153 \$10366 \$9059 \$10112 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34661 \$16 \$10446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34662 \$153 \$10425 \$10397 \$10446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34664 \$16 \$10467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34665 \$153 \$10452 \$10397 \$10467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34666 \$153 \$10426 \$10397 \$10392 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34667 \$153 \$9713 \$8977 \$9646 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34668 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$34670 \$16 \$10392 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34671 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$34673 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$34674 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$34675 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$34676 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$34677 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$34678 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$34680 \$153 \$5990 \$5896 \$5181 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34681 \$153 \$5917 \$5896 \$5403 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34682 \$16 \$5181 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34683 \$153 \$5768 \$5710 \$5736 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34685 \$16 \$5245 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34688 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$34689 \$153 \$5991 \$5896 \$5518 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34690 \$16 \$5736 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34692 \$153 \$5896 \$5376 \$5943 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$34693 \$16 \$4320 \$6051 \$5943 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$34694 \$16 \$5518 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34696 \$153 \$5975 \$4706 \$5837 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34697 \$153 \$5836 \$5373 \$5762 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34698 \$153 \$5991 \$5463 \$5837 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34700 \$153 \$5918 \$5710 \$5518 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34701 \$16 \$4742 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34702 \$153 \$5918 \$5463 \$5762 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34703 \$153 \$5790 \$5463 \$5618 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34705 \$153 \$5944 \$5976 \$5518 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34706 \$153 \$5870 \$5628 \$5736 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34707 \$153 \$5992 \$5055 \$5977 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34708 \$16 \$5489 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34709 \$16 \$5736 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34711 \$153 \$5945 \$5976 \$5245 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34714 \$153 \$5870 \$5055 \$5618 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34715 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$34716 \$153 \$5838 \$5107 \$5618 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34717 \$153 \$5945 \$5107 \$5977 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34718 \$153 \$5976 \$4269 \$5871 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$34719 \$16 \$4178 \$16 \$153 \$5977 VNB sky130_fd_sc_hd__inv_1
X$34720 \$16 \$5245 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34722 \$153 \$5732 \$5463 \$5619 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34723 \$153 \$6053 \$4616 \$5897 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$34724 \$153 \$6026 \$4706 \$6043 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34726 \$153 \$5946 \$6053 \$5403 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34727 \$16 \$4479 \$5712 \$5897 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$34730 \$153 \$5919 \$6053 \$5736 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34731 \$153 \$5946 \$5405 \$6043 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34732 \$16 \$5403 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34733 \$16 \$5736 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34735 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$34736 \$153 \$5978 \$5174 \$5993 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34737 \$153 \$6056 \$5388 \$5898 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$34739 \$16 \$4421 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34740 \$16 \$4421 \$5712 \$5898 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$34741 \$153 \$5920 \$5711 \$5736 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34742 \$153 \$5947 \$6056 \$5403 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34743 \$153 \$5994 \$4706 \$5993 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34744 \$16 \$5404 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34745 \$16 \$5736 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34748 \$153 \$5872 \$5711 \$5518 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34749 \$16 \$5403 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34750 \$16 \$4421 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34752 \$153 \$5995 \$5948 \$5403 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34753 \$153 \$5872 \$5463 \$5721 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34754 \$16 \$5404 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34755 \$153 \$5874 \$5349 \$5873 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$34758 \$153 \$5948 \$5230 \$5839 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$34759 \$153 \$5771 \$5645 \$5736 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34760 \$16 \$5403 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34761 \$153 \$5921 \$5874 \$5274 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34763 \$16 \$5736 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34765 \$153 \$5921 \$4706 \$5890 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34766 \$16 \$5274 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34768 \$153 \$5899 \$5874 \$5245 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34769 \$16 \$3198 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34770 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$34771 \$153 \$5899 \$5107 \$5890 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34772 \$16 \$4146 \$16 \$153 \$5890 VNB sky130_fd_sc_hd__inv_1
X$34773 \$16 \$5274 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34774 \$153 \$5875 \$5645 \$5274 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34776 \$153 \$5949 \$5645 \$5245 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34777 \$153 \$5875 \$4706 \$5621 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34778 \$153 \$6120 \$5228 \$5996 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$34779 \$16 \$5245 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34780 \$16 \$4869 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34782 \$16 \$5228 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34784 \$153 \$5832 \$4631 \$5792 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$34785 \$153 \$5979 \$5463 \$5722 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34786 \$153 \$5950 \$5832 \$5274 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34788 \$153 \$5922 \$5832 \$5404 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34790 \$16 \$5245 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34791 \$16 \$5489 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34792 \$153 \$5923 \$5832 \$5489 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34793 \$153 \$5922 \$5177 \$5722 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34794 \$16 \$5404 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34796 \$16 \$5181 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34797 \$153 \$5951 \$5832 \$5181 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34798 \$16 \$5403 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34800 \$16 \$4712 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34801 \$16 \$4320 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34803 \$153 \$5924 \$5832 \$5736 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34804 \$153 \$5951 \$5174 \$5722 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34805 \$153 \$5840 \$5405 \$5722 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34806 \$16 \$4320 \$5900 \$5841 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$34807 \$16 \$5736 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34809 \$153 \$5876 \$5833 \$5467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34810 \$16 \$5900 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34813 \$153 \$5952 \$5833 \$5271 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34814 \$16 \$5467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34815 \$16 \$5338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34816 \$153 \$5842 \$5209 \$5877 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34817 \$153 \$5952 \$5069 \$5877 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34818 \$16 \$4320 \$16 \$153 \$5877 VNB sky130_fd_sc_hd__inv_1
X$34819 \$16 \$5271 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34820 \$16 \$4742 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34822 \$16 \$4320 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34825 \$153 \$5953 \$5833 \$5469 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34826 \$153 \$5668 \$5287 \$5564 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34827 \$153 \$5699 \$5287 \$5622 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34828 \$153 \$5997 \$5205 \$5877 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34829 \$153 \$5843 \$5390 \$5877 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34831 \$16 \$5469 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34832 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$34834 \$153 \$5954 \$5901 \$5338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34835 \$153 \$5844 \$5901 \$5324 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34836 \$153 \$5998 \$5205 \$5845 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34837 \$16 \$5324 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34838 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$34841 \$16 \$4179 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34842 \$153 \$5954 \$5209 \$5845 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34844 \$153 \$5925 \$5901 \$5271 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34845 \$153 \$5968 \$5287 \$5845 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34846 \$153 \$5999 \$5406 \$5845 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34847 \$153 \$5925 \$5069 \$5845 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34849 \$16 \$4616 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34850 \$16 \$5271 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34851 \$16 \$4229 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34853 \$153 \$5955 \$5669 \$5478 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34854 \$153 \$5926 \$5669 \$5232 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34855 \$153 \$5926 \$5205 \$5623 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34856 \$16 \$4479 \$5713 \$5847 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$34857 \$16 \$5232 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34859 \$153 \$5927 \$5669 \$5469 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34860 \$153 \$5956 \$5669 \$5467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34861 \$153 \$5956 \$5406 \$5623 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34862 \$153 \$5927 \$5287 \$5623 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34863 \$16 \$5467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34864 \$16 \$5469 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34865 \$16 \$5388 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34869 \$153 \$5928 \$5653 \$5566 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34870 \$153 \$5957 \$5849 \$5271 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34871 \$153 \$5850 \$5390 \$5595 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34872 \$153 \$6000 \$5096 \$5980 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34873 \$16 \$5566 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34875 \$16 \$4421 \$16 \$153 \$5980 VNB sky130_fd_sc_hd__inv_1
X$34876 \$153 \$5928 \$5519 \$5595 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34877 \$16 \$5271 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34879 \$16 \$4600 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34880 \$16 \$5230 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34881 \$16 \$4600 \$5713 \$5969 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$34883 \$153 \$5851 \$5205 \$5595 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34884 \$153 \$6001 \$5230 \$5969 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$34885 \$16 \$5349 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34886 \$153 \$5929 \$5349 \$5958 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$34888 \$16 \$4146 \$5713 \$5958 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$34890 \$153 \$5829 \$5929 \$5324 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34891 \$153 \$5828 \$5929 \$5467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34893 \$16 \$3064 \$16 \$153 \$5772 VNB sky130_fd_sc_hd__clkbuf_2
X$34894 \$153 \$5981 \$5069 \$5852 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34897 \$16 \$4146 \$16 \$153 \$5852 VNB sky130_fd_sc_hd__inv_1
X$34898 \$16 \$5324 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34899 \$16 \$5467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34901 \$153 \$5902 \$5673 \$5566 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34902 \$153 \$5930 \$5673 \$5478 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34903 \$16 \$5566 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34904 \$16 \$5478 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34905 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$34906 \$153 \$5853 \$5406 \$5726 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34908 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$34910 \$153 \$5902 \$5519 \$5726 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34911 \$153 \$6002 \$5390 \$5982 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34912 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$34913 \$153 \$5983 \$5069 \$5982 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34914 \$16 \$5065 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34915 \$153 \$5854 \$5287 \$5631 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34917 \$153 \$5984 \$5406 \$5982 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34919 \$16 \$5324 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34920 \$16 \$5469 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34921 \$16 \$5228 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34922 \$153 \$5830 \$5065 \$5970 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$34923 \$153 \$5878 \$5549 \$5566 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34924 \$16 \$4712 \$5479 \$5970 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$34926 \$153 \$5774 \$5830 \$5566 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34927 \$16 \$5566 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34928 \$16 \$5478 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34930 \$153 \$6003 \$5830 \$5478 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34932 \$153 \$5855 \$5205 \$5815 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34933 \$16 \$5467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34934 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$34935 \$16 \$5566 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34936 \$153 \$5959 \$5830 \$5271 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34937 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$34938 \$16 \$5469 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34940 \$153 \$5931 \$5830 \$5469 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34941 \$153 \$5959 \$5069 \$5815 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34942 \$153 \$5931 \$5287 \$5815 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34943 \$153 \$6004 \$5096 \$5815 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34945 \$153 \$5879 \$5632 \$5796 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34948 \$153 \$5903 \$6067 \$5605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34949 \$153 \$5903 \$5625 \$6005 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34950 \$16 \$5605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34951 \$16 \$5714 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34953 \$16 \$5856 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34954 \$16 \$5932 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34955 \$153 \$5960 \$6067 \$5856 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34957 \$16 \$5856 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34959 \$153 \$5933 \$5632 \$5856 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34960 \$153 \$5960 \$5795 \$6005 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34961 \$16 \$5528 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34962 \$153 \$5880 \$6067 \$5528 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34963 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$34964 \$16 \$5702 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34966 \$153 \$5904 \$6067 \$5702 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34967 \$153 \$5880 \$5500 \$6005 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34968 \$153 \$5904 \$5470 \$6005 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34969 \$153 \$6067 \$4430 \$5971 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$34970 \$16 \$4324 \$16 \$153 \$6005 VNB sky130_fd_sc_hd__inv_1
X$34973 \$16 \$4324 \$5428 \$5971 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$34974 \$16 \$5819 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34975 \$153 \$6006 \$5961 \$5819 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34977 \$16 \$5834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34978 \$153 \$5857 \$6200 \$5340 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34979 \$153 \$5858 \$5881 \$5340 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34980 \$16 \$4430 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34981 \$16 \$4324 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34982 \$16 \$5856 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34983 \$153 \$5778 \$5655 \$5856 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34984 \$16 \$5702 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34986 \$153 \$5905 \$5961 \$5702 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$34987 \$153 \$5905 \$5470 \$5891 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34988 \$16 \$5834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34989 \$153 \$5961 \$4560 \$5934 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$34990 \$16 \$4432 \$5428 \$5934 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$34992 \$16 \$4432 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34993 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$34994 \$16 \$4432 \$16 \$153 \$5891 VNB sky130_fd_sc_hd__inv_1
X$34995 \$153 \$5859 \$5881 \$5571 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$34996 \$16 \$4560 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$34997 \$16 \$4415 \$5428 \$5972 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$34998 \$153 \$5973 \$4542 \$5972 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$34999 \$16 \$4432 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35000 \$16 \$4415 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35001 \$16 \$5834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35002 \$153 \$5882 \$5552 \$5834 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35004 \$153 \$6007 \$5755 \$6089 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35005 \$153 \$5860 \$6200 \$5472 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35007 \$153 \$6008 \$5973 \$5702 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35008 \$153 \$5882 \$5881 \$5472 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35012 \$153 \$5861 \$5795 \$5472 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35013 \$16 \$4415 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35014 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$35015 \$16 \$5796 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35016 \$153 \$6009 \$6011 \$5856 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35017 \$153 \$5781 \$5633 \$5796 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35018 \$16 \$5353 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35019 \$16 \$5856 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35020 \$153 \$5818 \$5881 \$5624 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35021 \$16 \$5714 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35023 \$153 \$6010 \$6011 \$5714 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35024 \$153 \$5797 \$5795 \$5624 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35025 \$16 \$4258 \$5906 \$5935 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$35026 \$153 \$6011 \$5264 \$5935 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$35027 \$16 \$5906 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35029 \$16 \$5834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35030 \$16 \$5796 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35032 \$153 \$5883 \$5656 \$5796 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35033 \$16 \$4258 \$16 \$153 \$5985 VNB sky130_fd_sc_hd__inv_1
X$35034 \$16 \$5605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35036 \$153 \$5986 \$5625 \$5985 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35037 \$153 \$5883 \$5775 \$5727 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35038 \$16 \$5264 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35039 \$16 \$4258 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35040 \$16 \$5906 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35041 \$16 \$4464 \$5906 \$5974 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$35042 \$153 \$5798 \$5795 \$5727 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35044 \$16 \$4464 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35045 \$153 \$6012 \$5381 \$5974 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$35046 \$153 \$5862 \$6200 \$5727 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35047 \$153 \$5884 \$5755 \$5892 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35049 \$153 \$6013 \$5658 \$5856 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35050 \$16 \$5856 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35051 \$16 \$5381 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35053 \$16 \$4464 \$16 \$153 \$5892 VNB sky130_fd_sc_hd__inv_1
X$35054 \$16 \$4464 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35055 \$153 \$5863 \$5881 \$5434 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35057 \$16 \$5796 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35058 \$153 \$5783 \$5658 \$5796 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35059 \$153 \$6013 \$5795 \$5434 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35061 \$16 \$5158 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35062 \$16 \$4724 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35063 \$16 \$5354 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35064 \$16 \$5906 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35065 \$16 \$5834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35067 \$16 \$5605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35068 \$153 \$5885 \$5634 \$5834 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35070 \$153 \$6014 \$5881 \$5987 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35071 \$16 \$5702 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35072 \$16 \$4376 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35073 \$16 \$5714 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35074 \$153 \$5885 \$5881 \$5574 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35075 \$16 \$4376 \$5906 \$6015 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$35076 \$153 \$5988 \$5470 \$5987 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35080 \$16 \$5528 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35082 \$153 \$5784 \$5634 \$5714 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35083 \$16 \$5796 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35084 \$153 \$6016 \$6072 \$5796 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35085 \$153 \$5864 \$5775 \$5574 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35086 \$16 \$4376 \$16 \$153 \$5987 VNB sky130_fd_sc_hd__inv_1
X$35088 \$16 \$5767 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35091 \$16 \$5636 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35092 \$153 \$5886 \$5907 \$5636 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35093 \$153 \$6017 \$5907 \$5767 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35094 \$153 \$5886 \$5509 \$5823 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35095 \$16 \$4430 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35096 \$153 \$5907 \$4430 \$5936 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$35099 \$16 \$4324 \$5485 \$5936 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$35100 \$16 \$5609 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35101 \$153 \$5962 \$5907 \$5609 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35102 \$153 \$5937 \$5907 \$5786 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35103 \$16 \$4093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35104 \$16 \$5786 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35105 \$16 \$5098 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35106 \$16 \$5786 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35107 \$16 \$4954 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35108 \$153 \$5708 \$5576 \$5786 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35110 \$153 \$5937 \$5635 \$5823 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35111 \$16 \$4780 \$16 \$153 \$6018 VNB sky130_fd_sc_hd__inv_1
X$35112 \$16 \$4780 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35113 \$16 \$4954 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35114 \$16 \$5767 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35115 \$16 \$3870 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35116 \$153 \$5909 \$5717 \$5767 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35117 \$153 \$5908 \$5806 \$5475 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35119 \$153 \$5909 \$5575 \$5475 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35120 \$153 \$5908 \$5717 \$5963 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35121 \$153 \$5939 \$5717 \$5887 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35122 \$16 \$5963 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35123 \$16 \$5786 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35124 \$16 \$5718 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35125 \$16 \$5887 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35126 \$16 \$1485 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35127 \$16 \$5887 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35129 \$153 \$5612 \$5074 \$5611 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35130 \$153 \$6019 \$5717 \$5718 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35131 \$153 \$5686 \$5938 \$5611 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35132 \$16 \$5887 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35134 \$153 \$5687 \$5806 \$5611 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35135 \$153 \$5835 \$4560 \$5940 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$35137 \$16 \$4432 \$5485 \$5940 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$35140 \$16 \$5963 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35141 \$16 \$5609 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35142 \$153 \$5888 \$5835 \$5963 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35143 \$16 \$5718 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35144 \$153 \$5964 \$5835 \$5718 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35145 \$16 \$4432 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35146 \$16 \$4432 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35147 \$153 \$5888 \$5806 \$5867 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35149 \$153 \$5964 \$5938 \$5867 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35150 \$16 \$5887 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35151 \$16 \$5579 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35153 \$153 \$5889 \$5835 \$5579 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35154 \$153 \$5965 \$5835 \$5887 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35156 \$153 \$5965 \$5627 \$5867 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35158 \$153 \$5889 \$5484 \$5867 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35159 \$153 \$5690 \$5627 \$5614 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35161 \$153 \$5910 \$5264 \$5911 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$35163 \$153 \$5868 \$5938 \$5559 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35164 \$16 \$4258 \$5582 \$5911 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$35165 \$16 \$5636 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35168 \$16 \$4258 \$16 \$153 \$5893 VNB sky130_fd_sc_hd__inv_1
X$35169 \$153 \$5912 \$5484 \$5893 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35170 \$153 \$6020 \$5910 \$5636 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35171 \$16 \$4258 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35173 \$153 \$5941 \$5381 \$5913 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$35174 \$16 \$4464 \$5582 \$5913 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$35176 \$16 \$5718 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35178 \$153 \$5966 \$5941 \$5718 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35179 \$153 \$5942 \$5941 \$5786 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35180 \$153 \$5942 \$5635 \$5894 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35181 \$153 \$5966 \$5938 \$5894 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35182 \$16 \$5887 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35183 \$153 \$4924 \$3719 \$3567 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35184 \$16 \$5579 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35186 \$153 \$6021 \$5941 \$5579 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35187 \$16 \$4316 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35188 \$16 \$5718 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35189 \$153 \$5914 \$5627 \$5894 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35190 \$153 \$6023 \$4316 \$6022 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$35191 \$153 \$5915 \$5575 \$5692 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35193 \$153 \$5915 \$5617 \$5767 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35194 \$16 \$5767 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35195 \$16 \$5718 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35196 \$153 \$5916 \$6023 \$5718 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35197 \$16 \$5718 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35199 \$153 \$5916 \$5938 \$5895 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35200 \$16 \$4376 \$16 \$153 \$5895 VNB sky130_fd_sc_hd__inv_1
X$35201 \$16 \$4376 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35206 \$16 \$5636 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35207 \$16 \$5786 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35208 \$153 \$5967 \$5617 \$5786 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35209 \$153 \$5869 \$5617 \$5636 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35211 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$35212 \$153 \$5989 \$5627 \$5895 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35214 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$35215 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$35217 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$35218 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$35219 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$35220 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$35221 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$35223 \$153 \$4382 \$4469 \$3616 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35224 \$153 \$4545 \$4469 \$3474 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35225 \$16 \$3616 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35226 \$16 \$3474 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35227 \$153 \$4545 \$3490 \$4372 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35228 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$35230 \$153 \$4629 \$3606 \$4372 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35232 \$153 \$4576 \$4469 \$3473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35233 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$35234 \$153 \$4649 \$4469 \$3571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35235 \$16 \$4320 \$4538 \$4486 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$35236 \$16 \$3473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35240 \$153 \$4487 \$3307 \$4372 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35241 \$16 \$3571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35242 \$16 \$4320 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35243 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$35244 \$16 \$3615 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35245 \$153 \$4650 \$4383 \$3615 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35246 \$16 \$4538 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35247 \$153 \$4577 \$4383 \$3474 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35249 \$153 \$4577 \$3490 \$4489 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35250 \$153 \$4578 \$4383 \$3473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35251 \$153 \$4578 \$3540 \$4489 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35253 \$153 \$4651 \$4614 \$3474 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35254 \$153 \$4418 \$3389 \$4489 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35256 \$153 \$4488 \$3478 \$4489 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35257 \$153 \$4653 \$4614 \$3473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35258 \$16 \$3474 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35260 \$16 \$4579 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35261 \$153 \$4471 \$4383 \$3709 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35263 \$16 \$4479 \$4144 \$4615 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$35266 \$153 \$4383 \$4616 \$4615 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$35267 \$153 \$4384 \$4383 \$3571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35268 \$16 \$4616 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35269 \$153 \$4547 \$4617 \$3616 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35270 \$153 \$4546 \$3307 \$4693 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35272 \$16 \$3571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35273 \$16 \$4479 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35275 \$153 \$4595 \$4617 \$3385 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35276 \$153 \$4547 \$3389 \$4527 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35277 \$153 \$4444 \$3490 \$4527 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35278 \$16 \$4621 \$4538 \$4654 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$35279 \$16 \$3474 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35280 \$153 \$4548 \$4617 \$3766 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35281 \$16 \$3385 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35283 \$153 \$4596 \$4617 \$3473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35284 \$153 \$4548 \$3478 \$4527 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35285 \$153 \$4596 \$3540 \$4527 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35286 \$16 \$3766 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35287 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$35288 \$16 \$3473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35290 \$16 \$3709 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35291 \$153 \$4387 \$4386 \$3473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35292 \$16 \$4538 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35293 \$16 \$4621 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35294 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$35296 \$153 \$4420 \$3389 \$4373 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35297 \$16 \$3473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35298 \$16 \$3474 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35299 \$153 \$4630 \$3394 \$4373 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35300 \$16 \$3616 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35302 \$153 \$4389 \$4386 \$3709 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35304 \$153 \$4656 \$4386 \$3615 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35305 \$153 \$4490 \$3478 \$4373 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35306 \$16 \$4600 \$4144 \$4657 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$35307 \$16 \$3709 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35308 \$16 \$3615 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35309 \$16 \$5230 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35310 \$153 \$4658 \$4390 \$3474 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35311 \$16 \$4600 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35314 \$153 \$4492 \$4390 \$3615 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35315 \$153 \$4491 \$3606 \$4329 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35316 \$16 \$3615 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35317 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$35318 \$16 \$3474 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35319 \$16 \$3385 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35320 \$16 \$3615 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35322 \$153 \$4493 \$4319 \$3615 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35323 \$16 \$3473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35325 \$153 \$4597 \$4390 \$3473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35326 \$153 \$4549 \$4319 \$3474 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35327 \$153 \$4597 \$3540 \$4329 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35329 \$16 \$4494 \$4012 \$4618 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$35331 \$153 \$4549 \$3490 \$4230 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35332 \$153 \$4319 \$4631 \$4618 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$35333 \$153 \$4422 \$3540 \$4230 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35334 \$16 \$3474 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35335 \$16 \$4494 \$16 \$153 \$4230 VNB sky130_fd_sc_hd__inv_1
X$35336 \$16 \$3473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35337 \$16 \$4528 \$16 \$153 \$4146 VNB sky130_fd_sc_hd__clkbuf_2
X$35338 \$16 \$5065 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35339 \$16 \$4712 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35340 \$16 \$4631 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35341 \$153 \$4528 \$4392 \$4447 \$4374 \$4393 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$35344 \$153 \$4619 \$4393 \$4447 \$4374 \$4392 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$35345 \$153 \$4495 \$4374 \$4447 \$4392 \$4393 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$35346 \$16 \$4550 \$16 \$153 \$4600 VNB sky130_fd_sc_hd__clkbuf_2
X$35347 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$35348 \$153 \$4374 \$4392 \$4550 \$4393 \$4447 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$35349 \$16 \$4447 \$4393 \$4374 \$4392 \$16 \$153 \$4660 VNB
+ sky130_fd_sc_hd__and4_2
X$35350 \$16 \$4037 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35351 \$16 \$4078 \$16 \$153 \$4393 VNB sky130_fd_sc_hd__clkbuf_2
X$35353 \$16 \$4184 \$16 \$153 \$4392 VNB sky130_fd_sc_hd__clkbuf_2
X$35355 \$16 \$4632 \$16 \$153 \$4447 VNB sky130_fd_sc_hd__clkbuf_2
X$35357 \$16 \$4496 \$4497 \$4539 \$153 \$16 \$4580 VNB sky130_fd_sc_hd__and3_4
X$35358 \$16 \$4580 \$16 \$153 \$4598 VNB sky130_fd_sc_hd__clkbuf_2
X$35359 \$16 \$4497 \$4539 \$4496 \$153 \$4632 \$16 VNB sky130_fd_sc_hd__and3b_4
X$35360 \$153 \$4497 \$4496 \$4581 \$4539 \$16 \$16 VNB sky130_fd_sc_hd__nor3b_4
X$35361 \$16 \$4620 \$16 \$153 \$4539 VNB sky130_fd_sc_hd__clkbuf_2
X$35362 \$16 \$4620 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35365 \$16 \$4161 \$16 \$153 \$3841 VNB sky130_fd_sc_hd__clkbuf_2
X$35366 \$16 \$4581 \$16 \$153 \$4662 VNB sky130_fd_sc_hd__clkbuf_2
X$35367 \$16 \$4812 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35368 \$16 \$4423 \$16 \$153 \$3638 VNB sky130_fd_sc_hd__clkbuf_2
X$35370 \$16 \$4621 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35372 \$153 \$4663 \$4540 \$3572 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35373 \$153 \$4582 \$4540 \$3621 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35374 \$16 \$3621 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35376 \$153 \$4582 \$3608 \$4633 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35378 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$35379 \$153 \$4583 \$4540 \$3573 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35380 \$16 \$4621 \$16 \$153 \$4633 VNB sky130_fd_sc_hd__inv_1
X$35381 \$16 \$4621 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35382 \$153 \$4551 \$4599 \$3480 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35383 \$16 \$3573 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35384 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$35386 \$153 \$4584 \$4599 \$3386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35388 \$153 \$4583 \$3079 \$4633 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35389 \$16 \$3480 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35390 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$35391 \$153 \$4664 \$4540 \$3386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35392 \$153 \$4551 \$3504 \$4529 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35393 \$16 \$3386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35394 \$16 \$4179 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35396 \$16 \$3386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35398 \$153 \$4522 \$4540 \$3492 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35399 \$153 \$4601 \$4540 \$3620 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35401 \$16 \$3620 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35402 \$153 \$4601 \$3645 \$4633 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35403 \$16 \$3480 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35405 \$153 \$4398 \$4616 \$4552 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$35407 \$16 \$4479 \$4014 \$4552 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$35408 \$16 \$4479 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35409 \$16 \$4479 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35410 \$16 \$3492 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35411 \$153 \$4554 \$4398 \$3480 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35412 \$16 \$4616 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35414 \$16 \$4479 \$16 \$153 \$4338 VNB sky130_fd_sc_hd__inv_1
X$35416 \$153 \$4553 \$3354 \$4338 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35417 \$153 \$4602 \$4398 \$3572 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35419 \$153 \$4554 \$3504 \$4338 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35420 \$16 \$3386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35421 \$153 \$4555 \$3556 \$4338 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35422 \$153 \$4602 \$3101 \$4338 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35423 \$16 \$4421 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35424 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$35425 \$16 \$3572 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35427 \$16 \$3621 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35430 \$153 \$4603 \$4622 \$3621 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35431 \$16 \$3543 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35432 \$153 \$4523 \$4322 \$3543 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35433 \$153 \$4604 \$4622 \$3620 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35434 \$153 \$4556 \$3079 \$4530 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35436 \$153 \$4339 \$4322 \$3480 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35437 \$153 \$4556 \$4622 \$3573 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35438 \$16 \$3480 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35439 \$16 \$4106 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35440 \$16 \$4600 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35441 \$16 \$4600 \$4014 \$4666 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$35443 \$153 \$4499 \$4541 \$3573 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35444 \$16 \$3573 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35447 \$153 \$4667 \$4541 \$3620 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35449 \$153 \$4585 \$4541 \$3621 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35450 \$16 \$4600 \$16 \$153 \$4498 VNB sky130_fd_sc_hd__inv_1
X$35451 \$16 \$3620 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35452 \$16 \$4600 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35454 \$153 \$4669 \$4541 \$3492 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35456 \$153 \$4586 \$4541 \$3543 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35457 \$153 \$4585 \$3608 \$4498 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35458 \$16 \$3621 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35459 \$16 \$3543 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35461 \$153 \$4480 \$4631 \$4557 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$35463 \$16 \$4494 \$3957 \$4557 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$35466 \$16 \$3492 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35467 \$16 \$4494 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35468 \$16 \$4494 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35469 \$153 \$4500 \$4480 \$3620 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35470 \$16 \$4631 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35472 \$153 \$4403 \$4480 \$3492 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35473 \$16 \$4494 \$16 \$153 \$4363 VNB sky130_fd_sc_hd__inv_1
X$35474 \$16 \$3492 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35475 \$16 \$3620 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35478 \$16 \$5228 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35479 \$153 \$4605 \$4480 \$3572 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35480 \$153 \$4341 \$4480 \$3573 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35481 \$153 \$4605 \$3101 \$4363 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35483 \$16 \$3621 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35484 \$16 \$3573 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35486 \$153 \$4524 \$4404 \$3573 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35487 \$16 \$3572 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35491 \$16 \$4869 \$16 \$153 \$4501 VNB sky130_fd_sc_hd__inv_1
X$35492 \$153 \$4672 \$4404 \$3621 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35493 \$153 \$4524 \$3079 \$4501 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35495 \$16 \$3621 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35496 \$153 \$4606 \$4404 \$3492 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35497 \$16 \$3572 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35498 \$16 \$3492 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35501 \$16 \$3573 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35503 \$153 \$4558 \$4404 \$3620 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35504 \$153 \$4606 \$3354 \$4501 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35505 \$153 \$4634 \$3645 \$4776 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35506 \$153 \$4558 \$3645 \$4501 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35510 \$16 \$3241 \$3310 \$3344 \$153 \$16 \$3983 VNB sky130_fd_sc_hd__and3_4
X$35511 \$153 \$4635 \$3556 \$4776 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35512 \$153 \$4559 \$3788 \$4531 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35513 \$153 \$4607 \$4481 \$4048 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35514 \$153 \$4429 \$3651 \$4531 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35516 \$153 \$4607 \$3858 \$4531 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35518 \$16 \$4048 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35519 \$153 \$4502 \$3716 \$4531 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35520 \$153 \$4457 \$3962 \$4531 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35521 \$16 \$3852 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35522 \$153 \$4503 \$4481 \$3852 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35523 \$16 \$3791 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35524 \$153 \$4673 \$3939 \$4531 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35526 \$16 \$3792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35527 \$16 \$3792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35528 \$16 \$4590 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35530 \$153 \$4481 \$4590 \$4674 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$35531 \$153 \$4504 \$3939 \$4234 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35532 \$153 \$4254 \$4430 \$4505 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$35533 \$153 \$4608 \$4722 \$3814 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35535 \$153 \$4431 \$4254 \$3731 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35536 \$153 \$4608 \$3651 \$4697 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35537 \$16 \$4048 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35538 \$153 \$4506 \$4165 \$4048 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35539 \$16 \$4675 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35540 \$16 \$3272 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35543 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$35544 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$35546 \$16 \$3852 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35547 \$16 \$4432 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35548 \$16 \$3731 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35549 \$153 \$4165 \$4560 \$4507 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$35550 \$16 \$4930 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35552 \$153 \$4623 \$3788 \$4587 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35553 \$153 \$4636 \$3788 \$4637 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35555 \$16 \$4432 \$16 \$153 \$4235 VNB sky130_fd_sc_hd__inv_1
X$35556 \$153 \$4508 \$3716 \$4235 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35557 \$153 \$4677 \$4698 \$4048 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35559 \$16 \$4475 \$16 \$153 \$4166 VNB sky130_fd_sc_hd__clkbuf_2
X$35560 \$153 \$4256 \$4542 \$4525 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$35561 \$16 \$3198 \$16 \$153 \$4475 VNB sky130_fd_sc_hd__clkbuf_2
X$35564 \$16 \$3198 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35565 \$16 \$3792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35567 \$153 \$4624 \$4638 \$3814 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35568 \$153 \$4561 \$4256 \$3792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35570 \$16 \$4542 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35571 \$16 \$4048 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35573 \$153 \$4678 \$4638 \$4048 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35574 \$16 \$4562 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35575 \$16 \$3889 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35577 \$153 \$4561 \$3939 \$4167 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35579 \$16 \$3791 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35580 \$153 \$4854 \$3716 \$4587 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35581 \$153 \$4588 \$4257 \$3889 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35582 \$153 \$4345 \$3651 \$4509 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35584 \$16 \$4562 \$16 \$153 \$4509 VNB sky130_fd_sc_hd__inv_1
X$35585 \$153 \$4588 \$3962 \$4509 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35586 \$153 \$4563 \$4257 \$3791 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35587 \$153 \$4280 \$3788 \$4509 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35588 \$153 \$4563 \$3919 \$4509 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35589 \$153 \$4624 \$3651 \$4587 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35591 \$153 \$4679 \$3919 \$4639 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35592 \$153 \$4564 \$4323 \$3792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35593 \$16 \$3792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35594 \$16 \$4609 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35596 \$16 \$4724 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35597 \$153 \$4564 \$3939 \$4236 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35598 \$16 \$3852 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35600 \$153 \$4640 \$3651 \$4639 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35602 \$153 \$4323 \$5381 \$4510 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$35604 \$16 \$4048 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35605 \$16 \$4464 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35607 \$16 \$3960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35608 \$153 \$4434 \$3788 \$4236 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35609 \$153 \$4566 \$4565 \$3889 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35610 \$153 \$4680 \$4565 \$3960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35612 \$16 \$3889 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35614 \$153 \$4566 \$3962 \$4532 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35615 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$35616 \$16 \$3852 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35617 \$153 \$4681 \$4565 \$3852 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35618 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$35619 \$16 \$4543 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35620 \$16 \$4567 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35621 \$16 \$3731 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35622 \$153 \$4526 \$4565 \$3731 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35623 \$16 \$4048 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35625 \$153 \$4682 \$4565 \$4048 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35626 \$153 \$4526 \$3788 \$4532 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35627 \$153 \$4683 \$4565 \$3791 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35628 \$16 \$3791 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35630 \$16 \$2233 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35631 \$16 \$4567 \$4015 \$4568 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$35633 \$153 \$4565 \$4784 \$4568 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$35634 \$153 \$4684 \$4565 \$3814 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35635 \$16 \$2387 \$16 \$153 \$4544 VNB sky130_fd_sc_hd__clkbuf_2
X$35636 \$153 \$4477 \$4544 \$4589 \$4436 \$16 \$16 VNB sky130_fd_sc_hd__nor3b_4
X$35637 \$16 \$4685 \$16 \$153 \$4324 VNB sky130_fd_sc_hd__clkbuf_2
X$35638 \$16 \$4305 \$16 \$153 \$4686 VNB sky130_fd_sc_hd__clkbuf_2
X$35640 \$16 \$4511 \$16 \$153 \$4610 VNB sky130_fd_sc_hd__clkbuf_2
X$35641 \$16 \$4625 \$16 \$153 \$4432 VNB sky130_fd_sc_hd__clkbuf_2
X$35642 \$16 \$4544 \$4477 \$4436 \$153 \$16 \$4569 VNB sky130_fd_sc_hd__and3_4
X$35643 \$153 \$4625 \$4730 \$4686 \$4641 \$4610 \$16 \$16 VNB
+ sky130_fd_sc_hd__nor4b_2
X$35644 \$16 \$3983 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35646 \$16 \$4348 \$16 \$153 \$4092 VNB sky130_fd_sc_hd__clkbuf_2
X$35647 \$16 \$5452 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35648 \$16 \$4512 \$16 \$153 \$4567 VNB sky130_fd_sc_hd__clkbuf_2
X$35649 \$153 \$4642 \$3565 \$3567 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35650 \$16 \$4930 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35653 \$16 \$4533 \$16 \$153 \$3929 VNB sky130_fd_sc_hd__clkbuf_2
X$35654 \$153 \$4611 \$4731 \$4057 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35655 \$153 \$4483 \$4590 \$4438 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$35656 \$16 \$4534 \$16 \$153 \$3870 VNB sky130_fd_sc_hd__clkbuf_2
X$35657 \$153 \$4687 \$3860 \$4643 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35659 \$16 \$3826 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35660 \$153 \$4535 \$4483 \$3721 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35662 \$16 \$4057 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35663 \$16 \$4057 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35664 \$16 \$4930 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35665 \$16 \$4057 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35666 \$153 \$4644 \$3719 \$4643 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35667 \$153 \$4535 \$3676 \$4378 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35668 \$16 \$4430 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35669 \$153 \$4612 \$4731 \$3721 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35670 \$16 \$3721 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35671 \$16 \$3898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35672 \$16 \$3602 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35674 \$153 \$4513 \$4731 \$3602 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35676 \$153 \$4645 \$3986 \$4643 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35677 \$16 \$3721 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35678 \$153 \$4612 \$3676 \$4643 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35680 \$16 \$3680 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35681 \$153 \$4570 \$4483 \$3680 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35682 \$16 \$4057 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35684 \$153 \$4571 \$4626 \$4057 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35685 \$153 \$4571 \$4414 \$4484 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35686 \$16 \$4613 \$16 \$153 \$3988 VNB sky130_fd_sc_hd__clkbuf_2
X$35687 \$153 \$4570 \$3719 \$4378 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35688 \$153 \$4325 \$4560 \$4514 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$35691 \$153 \$4572 \$4414 \$4369 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35692 \$16 \$3680 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35693 \$16 \$4129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35694 \$153 \$4350 \$4325 \$3680 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35695 \$153 \$4572 \$4325 \$4057 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35697 \$16 \$3691 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35698 \$153 \$4515 \$3142 \$4369 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35701 \$16 \$4057 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35702 \$16 \$3898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35703 \$153 \$4690 \$4627 \$4057 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35704 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$35705 \$16 \$3721 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35706 \$153 \$4536 \$4325 \$3721 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35707 \$153 \$4352 \$4325 \$3898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35710 \$153 \$4536 \$3676 \$4369 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35711 \$153 \$4267 \$4609 \$4691 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$35712 \$16 \$4613 \$16 \$153 \$4156 VNB sky130_fd_sc_hd__clkbuf_2
X$35714 \$153 \$4591 \$4267 \$4129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35715 \$16 \$4609 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35717 \$16 \$4129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35719 \$153 \$4128 \$3565 \$4379 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35720 \$16 \$4562 \$16 \$153 \$4857 VNB sky130_fd_sc_hd__inv_1
X$35722 \$153 \$4573 \$4267 \$3691 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35723 \$16 \$3691 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35725 \$16 \$5381 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35726 \$153 \$4268 \$5381 \$4628 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$35727 \$16 \$4464 \$4156 \$4628 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$35731 \$153 \$4647 \$3986 \$4646 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35732 \$16 \$4057 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35733 \$153 \$4592 \$4268 \$4057 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35734 \$153 \$4355 \$3565 \$4371 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35736 \$153 \$4131 \$3719 \$4371 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35737 \$153 \$4289 \$3986 \$4371 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35739 \$153 \$4518 \$3893 \$4371 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35740 \$153 \$4485 \$4784 \$4574 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$35741 \$153 \$4648 \$4414 \$4537 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35743 \$16 \$4129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35745 \$153 \$4575 \$3719 \$4537 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35746 \$153 \$4575 \$4485 \$3680 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35748 \$16 \$4567 \$4156 \$4574 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$35749 \$153 \$4519 \$3986 \$4537 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35750 \$16 \$4567 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35751 \$153 \$4468 \$3142 \$4537 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35752 \$153 \$4593 \$4485 \$3602 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35753 \$16 \$3602 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35754 \$153 \$4520 \$3893 \$4537 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35756 \$16 \$4057 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35757 \$16 \$3602 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35758 \$16 \$3721 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35759 \$16 \$3721 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35761 \$153 \$4594 \$4485 \$3721 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35762 \$153 \$4648 \$4485 \$4057 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35763 \$16 \$3898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35764 \$153 \$4357 \$3860 \$4173 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35765 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$35767 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$35768 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$35769 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$35770 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$35771 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$35772 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$35773 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$35774 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$35777 \$153 \$3776 \$3942 \$3616 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35778 \$153 \$4028 \$3942 \$3766 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35779 \$16 \$3474 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35780 \$153 \$3627 \$3708 \$3474 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35781 \$16 \$3766 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35784 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$35786 \$153 \$3944 \$3942 \$3473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35787 \$153 \$3943 \$3490 \$3765 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35788 \$16 \$3474 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35789 \$16 \$3616 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35790 \$16 \$3473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35791 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$35793 \$153 \$3993 \$3942 \$3571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35795 \$153 \$3944 \$3540 \$3765 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35797 \$16 \$3692 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35798 \$153 \$3993 \$3422 \$3765 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35800 \$153 \$3708 \$3660 \$3900 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$35801 \$16 \$3571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35802 \$16 \$3686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35803 \$16 \$4162 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35805 \$16 \$3571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35807 \$16 \$3638 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35808 \$16 \$3660 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35811 \$16 \$3686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35812 \$16 \$3638 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35813 \$153 \$3945 \$3864 \$3709 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35814 \$153 \$3994 \$3864 \$3571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35816 \$16 \$3571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35817 \$153 \$3994 \$3422 \$3934 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35818 \$16 \$3615 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35821 \$153 \$3945 \$3606 \$3934 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35823 \$153 \$3995 \$3864 \$3385 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35824 \$16 \$3709 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35825 \$153 \$3901 \$3864 \$3474 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35826 \$16 \$3473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35827 \$16 \$3385 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35828 \$16 \$4229 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35829 \$153 \$3901 \$3490 \$3934 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35831 \$153 \$3995 \$3394 \$3934 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35832 \$16 \$3474 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35833 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$35834 \$16 \$3778 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35835 \$153 \$3946 \$3845 \$3474 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35837 \$153 \$4029 \$3845 \$3766 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35840 \$153 \$3946 \$3490 \$3872 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35841 \$153 \$4030 \$3845 \$3615 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35842 \$16 \$3474 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35843 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$35844 \$16 \$3615 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35846 \$153 \$3969 \$3845 \$3709 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35847 \$153 \$4018 \$3540 \$3872 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35849 \$153 \$3969 \$3606 \$3872 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35850 \$16 \$3709 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35851 \$16 \$3686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35852 \$153 \$4031 \$3947 \$3474 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35853 \$16 \$3616 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35854 \$153 \$3902 \$3947 \$3709 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35855 \$16 \$3474 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35856 \$16 \$3709 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35858 \$153 \$3902 \$3606 \$3875 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35860 \$16 \$5095 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35862 \$153 \$3996 \$3947 \$3473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35863 \$153 \$3903 \$3947 \$3571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35864 \$16 \$3473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35866 \$16 \$3997 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35867 \$153 \$3769 \$3499 \$3709 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35868 \$16 \$3997 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35870 \$153 \$3996 \$3540 \$3875 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35871 \$153 \$4033 \$3838 \$3385 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35872 \$16 \$3709 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35873 \$16 \$3997 \$16 \$153 \$3409 VNB sky130_fd_sc_hd__inv_1
X$35875 \$153 \$3904 \$3307 \$3935 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35876 \$153 \$4035 \$3838 \$3709 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35878 \$153 \$3846 \$3422 \$3935 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35880 \$153 \$3410 \$3949 \$3948 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$35881 \$153 \$4035 \$3606 \$3935 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35882 \$16 \$3658 \$4012 \$3948 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$35883 \$153 \$3970 \$4077 \$3385 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35886 \$16 \$3949 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35888 \$16 \$3473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35889 \$153 \$3970 \$3394 \$4019 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35890 \$153 \$3172 \$1815 \$2743 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35891 \$153 \$4036 \$4077 \$3766 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35892 \$16 \$3385 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35893 \$16 \$3907 \$4012 \$3950 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$35896 \$16 \$3907 \$16 \$153 \$3607 VNB sky130_fd_sc_hd__inv_1
X$35897 \$153 \$3998 \$4077 \$3709 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35898 \$153 \$3725 \$3906 \$3950 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$35899 \$16 \$3709 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35900 \$153 \$3998 \$3606 \$4019 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35901 \$153 \$3908 \$3725 \$3709 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35904 \$16 \$3886 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35906 \$16 \$3615 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35907 \$16 \$16 \$153 VNB sky130_fd_sc_hd__conb_1
X$35908 \$153 \$3908 \$3606 \$3607 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35909 \$153 \$153 \$3422 \$4020 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35910 \$153 \$3951 \$3307 \$3607 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35911 \$153 \$153 \$3394 \$4020 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35912 \$16 \$3781 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35913 \$16 \$3866 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35915 \$16 \$3711 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35917 \$16 \$3867 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35918 \$16 \$3953 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35919 \$16 \$3726 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35920 \$16 \$3712 \$4037 \$3805 \$3837 \$16 \$153 VNB sky130_fd_sc_hd__mux2_1
X$35921 \$16 \$3712 \$3910 \$3909 \$713 \$16 \$153 VNB sky130_fd_sc_hd__mux2_1
X$35923 \$16 \$3418 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35924 \$16 \$2634 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35925 \$16 \$3418 \$16 \$153 \$3712 VNB sky130_fd_sc_hd__clkbuf_2
X$35926 \$153 \$3591 \$3971 \$3553 \$3952 \$3953 \$3770 \$3592 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$35927 \$16 \$3778 \$3783 \$4038 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$35928 \$16 \$3783 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35931 \$16 \$3712 \$4039 \$3971 \$233 \$16 \$153 VNB sky130_fd_sc_hd__mux2_1
X$35932 \$153 \$3972 \$3785 \$3572 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35933 \$16 \$3778 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35934 \$16 \$3770 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35935 \$16 \$3638 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35936 \$16 \$3778 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35937 \$16 \$3572 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35938 \$153 \$3876 \$3785 \$3573 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35939 \$16 \$3778 \$16 \$153 \$3868 VNB sky130_fd_sc_hd__inv_1
X$35941 \$153 \$3936 \$3785 \$3543 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35942 \$153 \$3972 \$3101 \$3868 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35943 \$153 \$3936 \$3556 \$3868 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35944 \$16 \$3543 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35945 \$153 \$4021 \$3079 \$4022 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35946 \$153 \$3973 \$3785 \$3620 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35949 \$153 \$3999 \$3785 \$3480 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35950 \$153 \$3973 \$3645 \$3868 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35951 \$153 \$3999 \$3504 \$3868 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35952 \$16 \$3620 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35953 \$16 \$3480 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35955 \$16 \$3910 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35956 \$153 \$3878 \$3954 \$3386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35958 \$153 \$3974 \$3954 \$3480 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35959 \$153 \$3974 \$3504 \$4068 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35960 \$16 \$3480 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35961 \$16 \$3841 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35963 \$153 \$3975 \$3954 \$3573 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35964 \$16 \$3386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35966 \$16 \$3543 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35968 \$153 \$4041 \$3954 \$3492 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35969 \$16 \$3573 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35970 \$16 \$5095 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35971 \$153 \$3413 \$5095 \$3912 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$35972 \$16 \$3492 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35973 \$153 \$4042 \$3955 \$3621 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35976 \$153 \$3938 \$3504 \$3937 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35977 \$153 \$3938 \$3955 \$3480 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35978 \$153 \$3976 \$3955 \$3386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35979 \$16 \$3879 \$3783 \$4013 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$35980 \$153 \$3850 \$3079 \$3937 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35983 \$153 \$3976 \$3435 \$3937 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35984 \$16 \$3386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35985 \$16 \$3714 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35986 \$153 \$3880 \$3869 \$3573 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35987 \$153 \$3977 \$3869 \$3620 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35988 \$153 \$3977 \$3645 \$3881 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$35991 \$16 \$3620 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35992 \$16 \$3573 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35993 \$16 \$3978 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35994 \$16 \$3543 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35995 \$16 \$1485 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$35997 \$153 \$3913 \$3869 \$3480 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35998 \$153 \$3882 \$3869 \$3386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$35999 \$153 \$3913 \$3504 \$3881 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36000 \$16 \$3386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36003 \$16 \$4146 \$4014 \$4043 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$36004 \$16 \$3480 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36005 \$16 \$4146 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36006 \$16 \$4146 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36008 \$153 \$3979 \$3956 \$3480 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36009 \$153 \$3883 \$3956 \$3386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36010 \$16 \$4146 \$16 \$153 \$3884 VNB sky130_fd_sc_hd__inv_1
X$36011 \$153 \$3979 \$3504 \$3884 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36013 \$16 \$3480 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36015 \$153 \$3980 \$3956 \$3543 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36016 \$16 \$3386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36017 \$153 \$3810 \$3556 \$3340 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36018 \$153 \$3980 \$3556 \$3884 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36019 \$16 \$3543 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36020 \$16 \$3658 \$3957 \$3885 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$36021 \$16 \$3621 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36023 \$153 \$3914 \$3956 \$3492 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36026 \$153 \$3887 \$3956 \$3573 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36027 \$153 \$3914 \$3354 \$3884 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36028 \$16 \$3573 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36029 \$16 \$3906 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36030 \$153 \$3787 \$3906 \$3981 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$36031 \$16 \$3492 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36034 \$16 \$3907 \$3957 \$3981 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$36035 \$16 \$3907 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36036 \$153 \$3584 \$3787 \$3386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36037 \$153 \$3915 \$3787 \$3572 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36038 \$16 \$3386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36039 \$153 \$3915 \$3101 \$3585 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36040 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$36042 \$153 \$3730 \$3787 \$3543 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36044 \$153 \$3982 \$3787 \$3621 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36045 \$16 \$3543 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36046 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$36047 \$16 \$3621 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36048 \$16 \$3272 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36050 \$16 \$3919 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36051 \$153 \$1539 \$3620 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$36052 \$16 \$3858 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36055 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36056 \$153 \$3866 \$1482 \$3716 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36057 \$153 \$3982 \$3608 \$3585 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36058 \$153 \$3953 \$1482 \$3858 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36059 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36060 \$16 \$1539 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36062 \$153 \$3096 \$3731 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$36063 \$153 \$3781 \$1482 \$1715 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36064 \$153 \$3634 \$1482 \$3763 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36065 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36067 \$16 \$3333 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36069 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36070 \$153 \$3555 \$1482 \$3788 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36071 \$153 \$4000 \$3958 \$3960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36072 \$16 \$2438 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36073 \$16 \$1558 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36074 \$16 \$1613 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36075 \$153 \$3917 \$3958 \$3791 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36076 \$16 \$4048 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36077 \$16 \$3852 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36079 \$153 \$4000 \$3716 \$3762 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36080 \$153 \$4118 \$3939 \$3762 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36081 \$153 \$3918 \$3958 \$3814 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36082 \$16 \$4093 \$16 \$153 \$3762 VNB sky130_fd_sc_hd__inv_1
X$36083 \$16 \$3960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36085 \$16 \$4048 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36086 \$153 \$4001 \$3715 \$4048 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36088 \$153 \$3918 \$3651 \$3762 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36089 \$16 \$3814 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36090 \$16 \$3791 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36091 \$153 \$3984 \$3715 \$3791 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36092 \$153 \$4001 \$3858 \$3160 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36093 \$16 \$3272 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36095 \$16 \$3792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36097 \$153 \$4314 \$3715 \$3889 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36098 \$153 \$3984 \$3919 \$3160 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36099 \$153 \$3959 \$3790 \$3792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36101 \$153 \$3816 \$3651 \$3890 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36103 \$16 \$3889 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36105 \$16 \$3960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36106 \$153 \$3959 \$3939 \$3890 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36107 \$153 \$4002 \$3790 \$3960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36108 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$36109 \$153 \$3817 \$3919 \$3890 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36110 \$153 \$4002 \$3716 \$3890 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36111 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$36112 \$16 \$3960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36113 \$153 \$3920 \$3622 \$3960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36117 \$16 \$3889 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36118 \$16 \$4047 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36119 \$16 \$4048 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36120 \$153 \$4003 \$3622 \$4048 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36121 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$36122 \$153 \$3920 \$3716 \$3732 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36123 \$153 \$4003 \$3858 \$3732 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36126 \$153 \$3961 \$3962 \$3732 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36128 \$16 \$3960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36129 \$153 \$4004 \$3717 \$3960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36130 \$16 \$3791 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36131 \$153 \$3921 \$3717 \$3791 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36132 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$36133 \$153 \$3921 \$3919 \$3773 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36135 \$153 \$4004 \$3716 \$3773 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36137 \$16 \$4048 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36139 \$153 \$3922 \$3670 \$4048 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36140 \$153 \$3963 \$3670 \$3791 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36142 \$16 \$3791 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36144 \$153 \$3857 \$3939 \$3891 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36145 \$153 \$3922 \$3858 \$3891 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36146 \$153 \$3963 \$3919 \$3891 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36147 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$36148 \$16 \$4016 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36149 \$16 \$4048 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36151 \$153 \$3923 \$3649 \$4048 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36152 \$16 \$4016 \$4015 \$4051 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$36153 \$16 \$3960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36154 \$16 \$3791 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36156 \$153 \$4005 \$3649 \$3791 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36157 \$153 \$3924 \$3649 \$3792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36158 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$36160 \$16 \$3960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36161 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$36162 \$153 \$3892 \$3718 \$3960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36163 \$16 \$3731 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36165 \$153 \$3924 \$3939 \$3609 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36166 \$16 \$3852 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36168 \$153 \$3985 \$4091 \$3852 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36169 \$153 \$4023 \$3716 \$4024 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36170 \$16 \$5002 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36171 \$16 \$3834 \$4015 \$4025 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$36172 \$16 \$4048 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36174 \$16 \$3559 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36175 \$153 \$3718 \$5002 \$4025 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$36176 \$153 \$3925 \$3718 \$4048 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36177 \$16 \$3791 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36179 \$16 \$3791 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36180 \$153 \$3925 \$3858 \$3610 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36181 \$153 \$4053 \$4091 \$3791 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36183 \$16 \$3834 \$16 \$153 \$3610 VNB sky130_fd_sc_hd__inv_1
X$36184 \$153 \$3940 \$3651 \$4024 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36185 \$153 \$3940 \$4091 \$3814 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36186 \$16 \$3086 \$3964 \$3673 \$3419 \$16 \$153 VNB sky130_fd_sc_hd__mux2_1
X$36187 \$16 \$3565 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36188 \$153 \$153 \$3565 \$3941 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36190 \$16 \$3983 \$16 \$153 \$3941 VNB sky130_fd_sc_hd__clkbuf_2
X$36192 \$153 \$153 \$3893 \$3941 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36193 \$16 \$3983 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36194 \$16 \$3834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36195 \$153 \$153 \$3719 \$3941 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36196 \$16 \$16 \$153 VNB sky130_fd_sc_hd__conb_1
X$36198 \$16 \$4026 \$16 \$153 \$3834 VNB sky130_fd_sc_hd__clkbuf_2
X$36199 \$16 \$3826 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36200 \$153 \$3795 \$4276 \$4054 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$36201 \$153 \$3926 \$3893 \$3461 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36203 \$16 \$3243 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36205 \$153 \$4006 \$3795 \$3826 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36206 \$153 \$3894 \$3795 \$3898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36207 \$153 \$4006 \$3893 \$3586 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36208 \$153 \$3927 \$3795 \$4057 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36210 \$153 \$3508 \$4129 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$36211 \$153 \$3987 \$3795 \$4129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36212 \$153 \$4027 \$3565 \$4072 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36213 \$16 \$4129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36214 \$16 \$3691 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36217 \$153 \$3705 \$4196 \$3966 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$36218 \$16 \$4057 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36220 \$153 \$4058 \$4017 \$3721 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36221 \$16 \$4139 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36222 \$16 \$3870 \$16 \$153 \$3461 VNB sky130_fd_sc_hd__inv_1
X$36223 \$16 \$3721 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36224 \$16 \$3721 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36225 \$153 \$3793 \$3705 \$3721 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36226 \$16 \$4196 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36227 \$16 \$3870 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36228 \$16 \$3898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36230 \$153 \$3896 \$4017 \$3898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36232 \$16 \$3898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36233 \$153 \$4154 \$3705 \$3898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36234 \$16 \$3929 \$3988 \$4007 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$36235 \$153 \$3796 \$4047 \$4007 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$36238 \$153 \$3755 \$3719 \$3775 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36240 \$16 \$4129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36241 \$153 \$3989 \$3796 \$4129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36242 \$153 \$3928 \$3676 \$3775 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36243 \$153 \$3989 \$3986 \$3775 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36244 \$16 \$3929 \$16 \$153 \$3775 VNB sky130_fd_sc_hd__inv_1
X$36248 \$16 \$3826 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36249 \$16 \$3898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36250 \$153 \$4061 \$3796 \$3898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36251 \$153 \$3990 \$3796 \$3826 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36253 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$36254 \$16 \$3826 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36255 \$153 \$4062 \$3623 \$3826 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36257 \$16 \$4057 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36258 \$16 \$3680 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36259 \$153 \$4073 \$3623 \$3680 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36260 \$153 \$3897 \$3623 \$4057 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36261 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$36262 \$153 \$3681 \$3565 \$3930 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36266 \$16 \$4258 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36267 \$16 \$3826 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36268 \$153 \$4008 \$3624 \$3826 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36269 \$153 \$3991 \$3624 \$3898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36270 \$153 \$4008 \$3893 \$3930 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36271 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$36274 \$153 \$3967 \$3986 \$3930 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36276 \$16 \$4016 \$4156 \$4063 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$36277 \$16 \$3826 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36278 \$153 \$3968 \$3722 \$3826 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36279 \$16 \$4016 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36280 \$153 \$3832 \$3719 \$3764 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36281 \$153 \$3968 \$3893 \$3764 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36282 \$16 \$4016 \$16 \$153 \$3764 VNB sky130_fd_sc_hd__inv_1
X$36284 \$153 \$4064 \$3722 \$3898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36286 \$16 \$3834 \$4156 \$3932 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$36287 \$153 \$3625 \$5002 \$3932 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$36288 \$153 \$3682 \$3565 \$3764 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36290 \$16 \$3602 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36292 \$16 \$4129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36293 \$153 \$4009 \$3871 \$3602 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36295 \$153 \$3933 \$3871 \$4129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36296 \$153 \$4009 \$3565 \$3899 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36297 \$153 \$3933 \$3986 \$3899 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36298 \$16 \$4092 \$16 \$153 \$3899 VNB sky130_fd_sc_hd__inv_1
X$36300 \$16 \$3721 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36301 \$153 \$3992 \$3871 \$3826 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36304 \$153 \$4065 \$3871 \$3898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36305 \$16 \$3898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36307 \$153 \$3471 \$1936 \$3328 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36308 \$153 \$3992 \$3893 \$3899 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36310 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$36312 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$36313 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$36314 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$36315 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$36316 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$36317 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$36318 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$36319 \$153 \$9382 \$9650 \$9129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36320 \$153 \$9649 \$9650 \$8715 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36321 \$16 \$8715 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36322 \$153 \$8826 \$9458 \$8580 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36323 \$16 \$9129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36326 \$153 \$9649 \$8638 \$9392 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36327 \$153 \$9600 \$8912 \$9392 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36329 \$153 \$9602 \$9650 \$9026 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36330 \$153 \$9763 \$8194 \$9392 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36331 \$153 \$9545 \$9650 \$8724 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36333 \$153 \$9601 \$8885 \$9392 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36334 \$153 \$9602 \$8726 \$9392 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36335 \$153 \$9650 \$7884 \$9715 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$36336 \$153 \$9582 \$9469 \$8580 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36338 \$153 \$9470 \$9469 \$8828 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36339 \$153 \$9582 \$8194 \$9270 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36340 \$16 \$8580 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36341 \$16 \$8828 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36343 \$16 \$8715 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36344 \$153 \$9603 \$8209 \$9583 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36345 \$153 \$9393 \$9469 \$8715 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36348 \$153 \$9604 \$8885 \$9583 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36349 \$153 \$9679 \$8194 \$9583 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36350 \$16 \$8003 \$16 \$153 \$9270 VNB sky130_fd_sc_hd__inv_1
X$36351 \$16 \$8724 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36352 \$16 \$8423 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36353 \$153 \$10184 \$8726 \$9583 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36354 \$153 \$9546 \$9543 \$8580 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36355 \$16 \$8003 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36358 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$36359 \$16 \$8580 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36360 \$153 \$9680 \$8885 \$9449 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36361 \$16 \$7922 \$9547 \$9474 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$36362 \$153 \$9637 \$9543 \$9129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36363 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$36364 \$16 \$8271 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36365 \$153 \$9637 \$8737 \$9449 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36368 \$153 \$9564 \$8726 \$9449 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36369 \$153 \$9681 \$8209 \$9449 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36370 \$16 \$8715 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36372 \$16 \$9129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36373 \$153 \$9605 \$9459 \$8715 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36374 \$153 \$9638 \$9459 \$8436 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36376 \$16 \$8297 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36377 \$153 \$9066 \$8726 \$7816 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36378 \$16 \$7816 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36380 \$16 \$8144 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36381 \$153 \$9651 \$9459 \$8580 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36382 \$153 \$9605 \$8638 \$9321 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36383 \$16 \$7816 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36385 \$16 \$7973 \$16 \$153 \$9321 VNB sky130_fd_sc_hd__inv_1
X$36386 \$153 \$9651 \$8194 \$9321 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36387 \$16 \$9129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36389 \$153 \$9508 \$8912 \$9321 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36390 \$16 \$8580 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36391 \$153 \$9652 \$9606 \$8580 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36392 \$16 \$7663 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36394 \$16 \$9414 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36395 \$153 \$9584 \$9606 \$8950 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36396 \$16 \$8580 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36397 \$16 \$8117 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36398 \$16 \$7973 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36400 \$153 \$9652 \$8194 \$9585 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36401 \$153 \$9584 \$8912 \$9585 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36403 \$153 \$9595 \$8209 \$9585 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36404 \$16 \$7992 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36405 \$16 \$8715 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36406 \$153 \$9653 \$9606 \$8715 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36408 \$16 \$8724 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36409 \$16 \$9129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36411 \$16 \$8828 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36413 \$153 \$9460 \$9334 \$8828 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36414 \$153 \$9653 \$8638 \$9585 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36416 \$153 \$9682 \$9673 \$8828 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36417 \$153 \$9673 \$6887 \$9607 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$36419 \$153 \$9683 \$9673 \$8715 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36420 \$16 \$8715 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36422 \$153 \$9608 \$9384 \$8828 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36423 \$153 \$9654 \$8457 \$9836 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36424 \$16 \$8828 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36425 \$16 \$8061 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36426 \$16 \$8169 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36427 \$153 \$9655 \$9673 \$9026 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36430 \$153 \$9566 \$8638 \$9396 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36431 \$153 \$9608 \$8885 \$9396 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36432 \$153 \$9682 \$8885 \$9567 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36434 \$153 \$9397 \$9384 \$8724 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36435 \$16 \$9026 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36436 \$16 \$7535 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36437 \$16 \$7655 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36439 \$153 \$9685 \$9673 \$8724 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36440 \$16 \$7535 \$16 \$153 \$9567 VNB sky130_fd_sc_hd__inv_1
X$36441 \$16 \$8724 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36442 \$16 \$9371 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36443 \$153 \$9609 \$7655 \$9568 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$36444 \$153 \$9684 \$8912 \$9567 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36445 \$16 \$8724 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36448 \$153 \$9656 \$9609 \$8816 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36449 \$153 \$9639 \$9609 \$8890 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36450 \$16 \$8816 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36452 \$153 \$9656 \$8804 \$9533 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36453 \$153 \$9549 \$9356 \$8647 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36454 \$16 \$8886 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36456 \$16 \$8001 \$16 \$153 \$9451 VNB sky130_fd_sc_hd__inv_1
X$36457 \$153 \$9611 \$9609 \$8898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36458 \$153 \$9639 \$8277 \$9533 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36459 \$153 \$9610 \$8614 \$9451 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36460 \$16 \$8898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36461 \$16 \$8001 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36462 \$16 \$10008 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36463 \$16 \$8001 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36464 \$153 \$9657 \$9609 \$8686 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36465 \$16 \$8686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36467 \$153 \$9611 \$8789 \$9533 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36468 \$153 \$9612 \$8818 \$9533 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36469 \$153 \$9657 \$8651 \$9533 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36470 \$153 \$9613 \$8610 \$9451 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36471 \$16 \$8686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36472 \$16 \$8139 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36473 \$16 \$8167 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36474 \$153 \$9206 \$9481 \$8890 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36476 \$153 \$9614 \$9481 \$8898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36477 \$16 \$8890 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36478 \$16 \$8898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36479 \$153 \$9614 \$8789 \$9186 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36480 \$153 \$9616 \$9481 \$8886 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36481 \$16 \$8728 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36483 \$16 \$8886 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36484 \$153 \$9484 \$8297 \$9615 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$36485 \$16 \$8144 \$9371 \$9615 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$36487 \$153 \$9617 \$9484 \$8816 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36488 \$153 \$9616 \$8727 \$9186 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36490 \$153 \$9617 \$8804 \$9373 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36492 \$16 \$8144 \$16 \$153 \$9373 VNB sky130_fd_sc_hd__inv_1
X$36493 \$16 \$8816 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36494 \$16 \$9371 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36495 \$153 \$9618 \$8818 \$9373 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36496 \$153 \$9658 \$9484 \$8898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36497 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$36498 \$153 \$9619 \$8727 \$9373 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36499 \$153 \$9658 \$8789 \$9373 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36501 \$16 \$7973 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36503 \$16 \$8117 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36504 \$16 \$8898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36505 \$153 \$9551 \$9487 \$8886 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36506 \$153 \$9686 \$9487 \$8898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36507 \$153 \$9374 \$8277 \$9111 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36508 \$16 \$8898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36509 \$16 \$8886 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36512 \$16 \$8728 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36513 \$153 \$9596 \$8818 \$9586 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36515 \$153 \$9687 \$9487 \$8816 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36516 \$16 \$8119 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36517 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$36518 \$153 \$9515 \$8277 \$9421 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36519 \$153 \$9686 \$8789 \$9488 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36521 \$153 \$9620 \$9463 \$8647 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36522 \$16 \$8816 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36524 \$153 \$9621 \$9463 \$8556 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36525 \$153 \$9640 \$9463 \$8728 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36526 \$153 \$9620 \$8614 \$9421 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36529 \$153 \$9688 \$8651 \$9421 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36530 \$153 \$9621 \$8610 \$9421 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36532 \$153 \$9622 \$9403 \$8890 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36533 \$16 \$8728 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36534 \$16 \$7887 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36535 \$16 \$6753 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36536 \$153 \$9622 \$8277 \$9452 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36538 \$153 \$9689 \$8789 \$9452 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36540 \$153 \$9570 \$8614 \$9452 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36542 \$153 \$9660 \$6887 \$9659 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$36543 \$16 \$6903 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36545 \$153 \$9571 \$8651 \$9452 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36546 \$153 \$9552 \$9424 \$8886 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36547 \$16 \$7535 \$9400 \$9659 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$36549 \$16 \$8728 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36550 \$153 \$9690 \$9660 \$8556 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36551 \$153 \$9512 \$8610 \$9488 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36552 \$153 \$9513 \$8818 \$9488 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36553 \$153 \$9551 \$8727 \$9488 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36555 \$153 \$9721 \$8277 \$9488 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36556 \$153 \$9490 \$8651 \$9300 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36557 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$36559 \$16 \$8890 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36560 \$153 \$9572 \$8614 \$9300 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36561 \$16 \$10042 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36562 \$153 \$10042 \$7082 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$36563 \$16 \$8614 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36564 \$16 \$8610 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36565 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$36567 \$16 \$8670 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36568 \$16 \$10501 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36569 \$16 \$9031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36570 \$153 \$9340 \$9404 \$9275 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36571 \$153 \$6920 \$8568 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$36572 \$16 \$9275 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36574 \$16 \$8568 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36576 \$153 \$8568 \$9188 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$36578 \$16 \$6920 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36579 \$16 \$8807 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36580 \$153 \$9624 \$9404 \$9188 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36581 \$153 \$9691 \$9174 \$9453 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36582 \$153 \$9623 \$9133 \$9453 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36585 \$16 \$8078 \$16 \$153 \$9625 VNB sky130_fd_sc_hd__clkbuf_2
X$36587 \$153 \$153 \$9133 \$9625 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36589 \$153 \$9187 \$9405 \$9031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36590 \$153 \$153 \$8676 \$9625 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36592 \$16 \$9045 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36593 \$16 \$9031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36594 \$153 \$9662 \$8676 \$9587 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36595 \$16 \$8807 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36596 \$16 \$9253 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36598 \$16 \$9275 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36599 \$153 \$9926 \$8917 \$9587 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36600 \$153 \$9692 \$9174 \$9587 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36601 \$153 \$9406 \$9405 \$9253 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36602 \$153 \$9693 \$9150 \$9723 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$36603 \$16 \$7839 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36604 \$16 \$9188 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36606 \$153 \$9694 \$9047 \$9587 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36607 \$16 \$9150 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36608 \$153 \$9626 \$8842 \$9587 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36609 \$16 \$8220 \$16 \$153 \$9587 VNB sky130_fd_sc_hd__inv_1
X$36610 \$153 \$9430 \$9081 \$9031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36611 \$16 \$9031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36613 \$16 \$9045 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36614 \$153 \$9663 \$9674 \$9045 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36616 \$153 \$9407 \$9081 \$9188 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36617 \$153 \$9663 \$9174 \$9695 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36618 \$153 \$9674 \$8250 \$9431 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$36620 \$153 \$9627 \$8917 \$9695 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36621 \$153 \$9544 \$8136 \$9628 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$36624 \$153 \$9696 \$8917 \$9465 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36625 \$153 \$9629 \$9544 \$9031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36626 \$153 \$9497 \$9544 \$8807 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36627 \$153 \$9664 \$9544 \$8936 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36630 \$153 \$9629 \$9133 \$9465 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36631 \$16 \$8807 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36632 \$16 \$8136 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36633 \$16 \$9253 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36634 \$153 \$9664 \$8842 \$9465 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36635 \$153 \$9641 \$9466 \$9253 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36636 \$16 \$7994 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36638 \$16 \$9642 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36641 \$16 \$9031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36643 \$153 \$9641 \$9252 \$9325 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36644 \$16 \$9275 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36645 \$16 \$9214 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36646 \$153 \$9630 \$9466 \$9214 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36647 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$36649 \$16 \$9642 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36650 \$153 \$9752 \$8285 \$9697 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$36651 \$16 \$8316 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36653 \$153 \$9573 \$9278 \$9325 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36654 \$153 \$9597 \$9433 \$9275 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36655 \$153 \$9630 \$9047 \$9325 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36656 \$16 \$8807 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36657 \$153 \$9597 \$9278 \$9521 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36658 \$16 \$8285 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36660 \$16 \$8316 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36661 \$16 \$9214 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36665 \$153 \$9665 \$9433 \$9214 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36666 \$153 \$9588 \$9433 \$8807 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36667 \$153 \$9575 \$9133 \$9521 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36668 \$153 \$9665 \$9047 \$9521 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36672 \$153 \$9666 \$9408 \$9275 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36673 \$153 \$9588 \$8676 \$9521 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36674 \$16 \$9275 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36676 \$153 \$9631 \$9133 \$9409 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36677 \$153 \$9666 \$9278 \$9409 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36678 \$153 \$9589 \$9408 \$9253 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36679 \$16 \$9253 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36680 \$16 \$9188 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36682 \$153 \$9667 \$9408 \$9188 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36683 \$153 \$9589 \$9252 \$9409 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36684 \$16 \$8265 \$9733 \$9698 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$36685 \$16 \$8359 \$9733 \$9576 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$36687 \$16 \$9214 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36689 \$16 \$9188 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36690 \$153 \$9668 \$9524 \$9253 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36691 \$16 \$9045 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36693 \$153 \$9598 \$9524 \$9188 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36694 \$153 \$9668 \$9252 \$9555 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36695 \$153 \$9598 \$8917 \$9555 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36696 \$16 \$9253 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36697 \$16 \$7431 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36698 \$16 \$7431 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36700 \$16 \$9275 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36701 \$16 \$8807 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36703 \$153 \$9556 \$9524 \$8807 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36704 \$153 \$9669 \$9524 \$9275 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36705 \$153 \$9669 \$9278 \$9555 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36706 \$153 \$9362 \$8676 \$9328 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36707 \$16 \$7386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36708 \$153 \$9699 \$9133 \$9555 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36711 \$153 \$9578 \$9122 \$9439 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36712 \$16 \$8078 \$16 \$153 \$9701 VNB sky130_fd_sc_hd__clkbuf_2
X$36713 \$153 \$9440 \$9467 \$8893 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36715 \$153 \$153 \$8923 \$9701 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36716 \$16 \$8078 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36718 \$16 \$8187 \$9675 \$9670 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$36719 \$16 \$8893 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36721 \$16 \$7839 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36722 \$153 \$9702 \$7839 \$9670 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$36724 \$153 \$9632 \$8923 \$9439 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36725 \$153 \$9590 \$9467 \$9154 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36727 \$153 \$9632 \$9467 \$8879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36729 \$153 \$9590 \$9103 \$9439 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36730 \$16 \$8879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36731 \$16 \$8187 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36733 \$153 \$9671 \$9702 \$8844 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36734 \$153 \$9579 \$8965 \$9439 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36735 \$153 \$9557 \$9441 \$8893 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36736 \$16 \$8844 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36737 \$16 \$8708 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36739 \$16 \$9134 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36740 \$16 \$9150 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36741 \$153 \$9676 \$9150 \$9599 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$36742 \$16 \$8220 \$9675 \$9599 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$36743 \$153 \$9363 \$8923 \$9329 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36744 \$153 \$9558 \$9676 \$8893 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36745 \$16 \$8893 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36746 \$16 \$8220 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36747 \$16 \$7076 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36748 \$16 \$8081 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36751 \$16 \$8220 \$16 \$153 \$9560 VNB sky130_fd_sc_hd__inv_1
X$36752 \$16 \$8220 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36753 \$16 \$9550 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36754 \$153 \$9633 \$8923 \$9560 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36755 \$16 \$9550 \$16 \$153 \$9191 VNB sky130_fd_sc_hd__clkbuf_2
X$36756 \$153 \$9634 \$9676 \$8927 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36757 \$16 \$8893 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36758 \$153 \$9634 \$9256 \$9560 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36759 \$153 \$9677 \$8136 \$9591 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$36761 \$16 \$8927 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36762 \$153 \$9703 \$8965 \$9560 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36763 \$16 \$7904 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36764 \$16 \$7904 \$9675 \$9591 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$36765 \$16 \$8044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36766 \$16 \$8927 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36767 \$16 \$7904 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36768 \$153 \$9704 \$9677 \$8927 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36769 \$153 \$9635 \$9122 \$9592 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36771 \$16 \$7904 \$16 \$153 \$9592 VNB sky130_fd_sc_hd__inv_1
X$36772 \$16 \$8044 \$16 \$153 \$9411 VNB sky130_fd_sc_hd__inv_1
X$36773 \$16 \$9154 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36775 \$16 \$8044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36776 \$153 \$9593 \$9468 \$9154 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36778 \$16 \$8844 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36779 \$153 \$9705 \$9677 \$8844 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36780 \$153 \$9593 \$9103 \$9411 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36782 \$16 \$8893 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36783 \$16 \$8879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36785 \$153 \$9594 \$9468 \$8879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36787 \$153 \$9672 \$9468 \$8893 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36788 \$16 \$8705 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36789 \$153 \$9672 \$8996 \$9411 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36790 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$36793 \$153 \$9594 \$8923 \$9411 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36794 \$16 \$8165 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36795 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$36796 \$16 \$8927 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36797 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$36798 \$153 \$9706 \$9726 \$8927 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36799 \$16 \$9154 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36800 \$153 \$9563 \$9364 \$9154 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36802 \$16 \$8879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36804 \$153 \$9527 \$9256 \$9280 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36805 \$153 \$9636 \$9364 \$8879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36806 \$153 \$9707 \$8996 \$9708 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36807 \$153 \$9636 \$8923 \$9280 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36809 \$16 \$8844 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36810 \$153 \$9709 \$9678 \$8844 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36813 \$16 \$8316 \$9562 \$9643 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$36814 \$16 \$8927 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36816 \$153 \$9644 \$9316 \$9134 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36818 \$153 \$8455 \$7639 \$8266 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36819 \$153 \$9644 \$9122 \$9239 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36820 \$153 \$9540 \$8996 \$9239 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36822 \$16 \$8359 \$9562 \$9580 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$36823 \$16 \$9134 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36825 \$153 \$9645 \$9581 \$9134 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36826 \$16 \$8893 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36827 \$153 \$9710 \$9581 \$8893 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36828 \$16 \$8359 \$16 \$153 \$9646 VNB sky130_fd_sc_hd__inv_1
X$36829 \$16 \$8265 \$9562 \$9711 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$36830 \$16 \$8927 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36832 \$16 \$8879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36833 \$153 \$9712 \$9581 \$8879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36834 \$153 \$9647 \$9581 \$8927 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36835 \$153 \$9446 \$9122 \$9366 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36837 \$153 \$9528 \$9256 \$9366 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36838 \$16 \$9035 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36841 \$16 \$9034 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36842 \$153 \$9713 \$9581 \$9035 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36843 \$153 \$9648 \$9391 \$9034 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36844 \$153 \$9714 \$9581 \$8844 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36845 \$153 \$9447 \$9103 \$9366 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36847 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$36848 \$16 \$8844 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36849 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$36850 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$36851 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$36852 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$36853 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$36854 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$36855 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$36856 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$36858 \$153 \$375 \$64 \$504 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36862 \$16 \$504 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36863 \$153 \$375 \$561 \$88 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36864 \$153 \$315 \$64 \$395 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36865 \$153 \$64 \$531 \$448 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$36867 \$153 \$449 \$511 \$249 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36869 \$153 \$376 \$64 \$419 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36870 \$153 \$376 \$349 \$88 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36871 \$153 \$278 \$65 \$263 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36872 \$16 \$249 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36873 \$16 \$503 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36875 \$16 \$585 \$503 \$450 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$36876 \$153 \$203 \$59 \$89 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36877 \$153 \$355 \$65 \$419 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36878 \$16 \$585 \$16 \$153 \$89 VNB sky130_fd_sc_hd__inv_1
X$36879 \$153 \$247 \$377 \$89 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36880 \$16 \$419 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36881 \$16 \$585 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36882 \$16 \$585 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36885 \$153 \$451 \$182 \$504 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36887 \$153 \$355 \$349 \$89 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36888 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$36889 \$153 \$429 \$394 \$89 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36890 \$153 \$378 \$182 \$395 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36891 \$16 \$419 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36892 \$16 \$504 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36894 \$153 \$378 \$394 \$94 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36895 \$153 \$316 \$182 \$263 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36896 \$16 \$395 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36897 \$16 \$537 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36898 \$16 \$430 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36899 \$16 \$263 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36900 \$153 \$453 \$66 \$249 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36901 \$153 \$316 \$234 \$94 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36903 \$153 \$317 \$66 \$419 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36904 \$16 \$249 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36906 \$16 \$454 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36907 \$153 \$379 \$234 \$270 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36908 \$16 \$419 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36910 \$153 \$379 \$67 \$263 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36911 \$153 \$401 \$394 \$270 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36913 \$153 \$401 \$67 \$395 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36914 \$153 \$129 \$30 \$270 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36916 \$16 \$395 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36917 \$16 \$249 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36918 \$16 \$263 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36919 \$153 \$345 \$234 \$98 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36920 \$16 \$323 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36921 \$153 \$402 \$68 \$395 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36923 \$153 \$345 \$68 \$263 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36925 \$153 \$402 \$394 \$98 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36926 \$153 \$281 \$377 \$98 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36927 \$16 \$395 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36928 \$16 \$280 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36929 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$36930 \$16 \$263 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36931 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$36933 \$153 \$456 \$190 \$419 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36934 \$153 \$318 \$190 \$249 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36935 \$153 \$357 \$190 \$395 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36936 \$153 \$318 \$377 \$100 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36938 \$153 \$357 \$394 \$100 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36939 \$16 \$380 \$16 \$153 \$100 VNB sky130_fd_sc_hd__inv_1
X$36940 \$16 \$419 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36941 \$16 \$395 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36942 \$16 \$249 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36944 \$16 \$380 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36945 \$153 \$457 \$69 \$395 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36947 \$16 \$356 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36948 \$153 \$183 \$69 \$184 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36950 \$153 \$282 \$377 \$101 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36951 \$16 \$356 \$16 \$153 \$101 VNB sky130_fd_sc_hd__inv_1
X$36952 \$16 \$184 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36953 \$16 \$395 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36954 \$153 \$458 \$349 \$101 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36956 \$153 \$381 \$70 \$263 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36957 \$153 \$283 \$70 \$419 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36959 \$153 \$250 \$234 \$101 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36960 \$16 \$419 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36961 \$16 \$504 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36962 \$153 \$319 \$70 \$504 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36963 \$153 \$459 \$70 \$395 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36964 \$153 \$319 \$561 \$172 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36965 \$16 \$504 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36967 \$16 \$351 \$16 \$153 \$172 VNB sky130_fd_sc_hd__inv_1
X$36968 \$153 \$460 \$71 \$504 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36970 \$153 \$888 \$71 \$419 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36971 \$153 \$431 \$234 \$432 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36972 \$16 \$419 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36974 \$16 \$395 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36976 \$153 \$382 \$71 \$395 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36978 \$16 \$588 \$16 \$153 \$173 VNB sky130_fd_sc_hd__inv_1
X$36979 \$153 \$433 \$394 \$432 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36980 \$153 \$72 \$531 \$286 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$36981 \$153 \$285 \$59 \$173 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36982 \$153 \$320 \$420 \$187 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36986 \$153 \$461 \$420 \$209 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36987 \$153 \$287 \$35 \$174 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$36988 \$16 \$585 \$16 \$153 \$271 VNB sky130_fd_sc_hd__inv_1
X$36989 \$16 \$209 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36990 \$16 \$264 \$16 \$153 \$174 VNB sky130_fd_sc_hd__inv_1
X$36991 \$16 \$358 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36992 \$153 \$462 \$420 \$358 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36993 \$16 \$264 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$36996 \$153 \$321 \$420 \$73 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36997 \$153 \$463 \$420 \$212 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$36998 \$153 \$322 \$72 \$212 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37000 \$16 \$73 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37001 \$16 \$212 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37002 \$153 \$322 \$347 \$174 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37003 \$153 \$434 \$104 \$271 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37004 \$16 \$60 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37006 \$153 \$464 \$74 \$209 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37007 \$16 \$212 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37009 \$16 \$279 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37011 \$153 \$350 \$74 \$293 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37012 \$153 \$465 \$74 \$187 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37013 \$16 \$212 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37014 \$16 \$293 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37015 \$16 \$187 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37016 \$16 \$209 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37017 \$153 \$106 \$185 \$293 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37019 \$16 \$279 \$507 \$466 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$37021 \$153 \$467 \$185 \$212 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37022 \$153 \$350 \$35 \$175 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37023 \$16 \$212 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37024 \$153 \$289 \$346 \$105 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37026 \$153 \$403 \$192 \$358 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37029 \$16 \$323 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37030 \$16 \$358 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37031 \$153 \$324 \$192 \$212 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37032 \$153 \$404 \$192 \$293 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37033 \$153 \$210 \$104 \$186 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37034 \$16 \$323 \$555 \$468 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$37036 \$16 \$209 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37037 \$16 \$212 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37038 \$16 \$187 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37040 \$16 \$293 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37042 \$153 \$470 \$24 \$187 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37043 \$153 \$291 \$347 \$325 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37044 \$16 \$323 \$16 \$153 \$325 VNB sky130_fd_sc_hd__inv_1
X$37045 \$153 \$471 \$24 \$358 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37048 \$16 \$323 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37049 \$153 \$292 \$346 \$325 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37050 \$16 \$358 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37052 \$153 \$396 \$53 \$293 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37054 \$153 \$326 \$53 \$212 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37056 \$153 \$405 \$53 \$358 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37057 \$153 \$383 \$53 \$187 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37058 \$153 \$405 \$253 \$176 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37059 \$153 \$326 \$347 \$176 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37060 \$153 \$396 \$35 \$176 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37063 \$153 \$384 \$193 \$209 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37064 \$16 \$380 \$16 \$153 \$20 VNB sky130_fd_sc_hd__inv_1
X$37066 \$153 \$406 \$193 \$358 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37067 \$153 \$327 \$193 \$293 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37068 \$16 \$358 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37070 \$153 \$406 \$253 \$20 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37071 \$153 \$385 \$194 \$212 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37072 \$153 \$327 \$35 \$20 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37074 \$16 \$293 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37075 \$16 \$351 \$16 \$153 \$188 VNB sky130_fd_sc_hd__inv_1
X$37076 \$153 \$473 \$194 \$293 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37077 \$16 \$212 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37078 \$16 \$351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37081 \$153 \$328 \$194 \$358 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37083 \$16 \$60 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37084 \$153 \$474 \$421 \$187 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37085 \$153 \$139 \$215 \$188 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37086 \$153 \$328 \$253 \$188 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37088 \$16 \$187 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37090 \$16 \$652 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37091 \$16 \$209 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37092 \$153 \$435 \$104 \$436 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37093 \$153 \$217 \$54 \$329 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37094 \$16 \$652 \$16 \$153 \$329 VNB sky130_fd_sc_hd__inv_1
X$37095 \$153 \$294 \$35 \$329 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37096 \$153 \$475 \$421 \$212 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37097 \$16 \$18 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37099 \$153 \$386 \$75 \$358 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37100 \$153 \$476 \$421 \$18 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37101 \$153 \$295 \$347 \$329 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37102 \$16 \$212 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37103 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$37104 \$153 \$359 \$76 \$424 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37107 \$153 \$477 \$422 \$424 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37108 \$153 \$296 \$389 \$352 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37109 \$16 \$424 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37110 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$37111 \$16 \$424 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37112 \$153 \$478 \$422 \$82 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37113 \$16 \$426 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37114 \$16 \$426 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37116 \$153 \$359 \$353 \$352 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37117 \$16 \$426 \$16 \$153 \$352 VNB sky130_fd_sc_hd__inv_1
X$37118 \$16 \$82 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37119 \$153 \$76 \$387 \$360 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$37120 \$16 \$426 \$397 \$360 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$37121 \$153 \$297 \$388 \$352 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37123 \$16 \$387 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37124 \$16 \$145 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37126 \$153 \$330 \$61 \$145 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37127 \$153 \$437 \$21 \$501 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37128 \$153 \$299 \$389 \$111 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37129 \$16 \$145 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37132 \$16 \$241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37134 \$153 \$409 \$407 \$145 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37135 \$153 \$331 \$61 \$241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37136 \$153 \$331 \$388 \$111 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37137 \$153 \$142 \$21 \$111 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37138 \$16 \$265 \$268 \$332 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$37139 \$16 \$438 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37141 \$153 \$61 \$423 \$332 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$37142 \$153 \$333 \$77 \$241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37144 \$16 \$273 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37145 \$153 \$361 \$77 \$273 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37146 \$153 \$333 \$388 \$113 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37148 \$16 \$268 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37149 \$153 \$361 \$389 \$113 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37151 \$16 \$397 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37152 \$16 \$424 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37153 \$16 \$273 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37154 \$16 \$145 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37155 \$153 \$362 \$78 \$424 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37157 \$16 \$354 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37158 \$16 \$82 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37159 \$153 \$197 \$78 \$82 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37161 \$153 \$482 \$78 \$241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37162 \$153 \$362 \$353 \$115 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37163 \$153 \$300 \$266 \$115 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37164 \$16 \$273 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37165 \$153 \$483 \$189 \$273 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37166 \$16 \$145 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37167 \$16 \$241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37169 \$153 \$334 \$189 \$145 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37170 \$153 \$484 \$189 \$241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37171 \$153 \$363 \$353 \$485 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37172 \$16 \$151 \$268 \$439 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$37174 \$16 \$145 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37176 \$153 \$274 \$267 \$145 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37178 \$153 \$486 \$267 \$424 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37179 \$153 \$364 \$388 \$177 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37180 \$16 \$424 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37181 \$153 \$267 \$116 \$410 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$37183 \$16 \$79 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37185 \$16 \$80 \$16 \$153 \$177 VNB sky130_fd_sc_hd__inv_1
X$37186 \$153 \$304 \$389 \$177 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37187 \$153 \$81 \$608 \$487 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$37188 \$153 \$335 \$81 \$79 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37190 \$153 \$335 \$112 \$117 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37193 \$153 \$365 \$81 \$273 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37194 \$16 \$241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37195 \$153 \$336 \$81 \$241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37197 \$153 \$440 \$112 \$771 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37198 \$153 \$365 \$389 \$117 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37199 \$16 \$82 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37202 \$153 \$411 \$425 \$82 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37203 \$153 \$337 \$62 \$424 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37205 \$153 \$337 \$353 \$120 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37206 \$153 \$411 \$44 \$348 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37207 \$16 \$441 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37208 \$16 \$258 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37209 \$16 \$258 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37211 \$153 \$489 \$559 \$348 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37212 \$16 \$369 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37213 \$16 \$276 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37214 \$16 \$276 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37215 \$16 \$241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37216 \$153 \$222 \$112 \$120 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37218 \$16 \$241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37219 \$153 \$412 \$425 \$241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37220 \$153 \$366 \$112 \$348 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37222 \$153 \$412 \$388 \$348 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37223 \$153 \$367 \$266 \$348 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37226 \$16 \$309 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37227 \$16 \$426 \$369 \$490 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$37228 \$16 \$446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37229 \$153 \$338 \$83 \$309 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37230 \$16 \$426 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37231 \$153 \$243 \$398 \$258 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37233 \$153 \$390 \$83 \$509 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37234 \$153 \$413 \$23 \$442 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37235 \$153 \$338 \$703 \$121 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37236 \$153 \$414 \$391 \$310 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37239 \$153 \$368 \$391 \$149 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37240 \$153 \$414 \$223 \$442 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37241 \$153 \$225 \$398 \$121 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37243 \$16 \$446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37244 \$16 \$509 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37245 \$16 \$399 \$16 \$153 \$258 VNB sky130_fd_sc_hd__inv_1
X$37247 \$16 \$309 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37249 \$153 \$400 \$84 \$446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37250 \$153 \$339 \$84 \$309 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37251 \$153 \$443 \$371 \$442 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37252 \$153 \$226 \$23 \$258 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37253 \$16 \$446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37255 \$153 \$415 \$85 \$446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37257 \$16 \$509 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37259 \$16 \$369 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37260 \$16 \$63 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37261 \$153 \$308 \$549 \$122 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37262 \$153 \$415 \$393 \$122 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37263 \$153 \$392 \$85 \$63 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37265 \$16 \$265 \$16 \$153 \$122 VNB sky130_fd_sc_hd__inv_1
X$37267 \$153 \$392 \$57 \$122 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37268 \$16 \$354 \$369 \$370 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$37269 \$16 \$310 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37270 \$16 \$309 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37271 \$153 \$275 \$227 \$309 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37273 \$153 \$492 \$427 \$149 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37276 \$16 \$354 \$16 \$153 \$124 VNB sky130_fd_sc_hd__inv_1
X$37277 \$16 \$438 \$16 \$153 \$502 VNB sky130_fd_sc_hd__inv_1
X$37279 \$16 \$509 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37280 \$16 \$446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37281 \$153 \$493 \$227 \$509 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37282 \$153 \$340 \$227 \$446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37283 \$16 \$178 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37284 \$153 \$311 \$549 \$124 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37285 \$16 \$438 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37287 \$16 \$428 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37289 \$153 \$340 \$393 \$124 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37290 \$16 \$258 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37291 \$16 \$446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37292 \$153 \$341 \$86 \$446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37294 \$16 \$509 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37295 \$16 \$151 \$428 \$495 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$37296 \$153 \$496 \$86 \$509 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37298 \$16 \$80 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37299 \$16 \$116 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37301 \$16 \$80 \$428 \$497 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$37302 \$153 \$444 \$703 \$179 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37304 \$153 \$372 \$371 \$179 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37305 \$153 \$750 \$703 \$445 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37306 \$153 \$342 \$87 \$63 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37308 \$153 \$372 \$87 \$509 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37309 \$153 \$373 \$393 \$179 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37311 \$153 \$313 \$549 \$179 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37312 \$153 \$229 \$223 \$179 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37313 \$16 \$446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37315 \$153 \$416 \$50 \$446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37316 \$16 \$309 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37317 \$16 \$723 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37318 \$153 \$374 \$371 \$126 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37319 \$153 \$314 \$703 \$126 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37320 \$153 \$416 \$393 \$126 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37322 \$16 \$509 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37324 \$16 \$63 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37325 \$16 \$309 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37326 \$153 \$343 \$277 \$63 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37328 \$153 \$417 \$277 \$309 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37330 \$153 \$343 \$57 \$181 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37332 \$153 \$417 \$703 \$181 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37333 \$16 \$615 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37335 \$16 \$276 \$16 \$153 \$181 VNB sky130_fd_sc_hd__inv_1
X$37337 \$16 \$178 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37338 \$153 \$418 \$277 \$178 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37339 \$16 \$276 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37340 \$16 \$306 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37341 \$16 \$310 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37342 \$153 \$344 \$277 \$310 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37343 \$153 \$418 \$549 \$181 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37344 \$153 \$344 \$223 \$181 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37347 \$153 \$447 \$393 \$181 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37348 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$37349 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$37350 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$37351 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$37352 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$37354 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$37356 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$37357 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$37358 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$37359 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$37360 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$37361 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$37362 \$153 \$2807 \$2643 \$2006 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37363 \$153 \$2845 \$2643 \$1687 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37364 \$16 \$2006 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37365 \$16 \$1687 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37366 \$153 \$2686 \$1547 \$2343 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37367 \$16 \$1980 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37370 \$153 \$2735 \$2009 \$2343 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37372 \$153 \$2808 \$2643 \$1795 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37374 \$153 \$2846 \$2643 \$2024 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37375 \$16 \$1942 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37376 \$16 \$1795 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37377 \$16 \$1390 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37378 \$153 \$2846 \$2210 \$2785 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37380 \$16 \$2024 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37381 \$153 \$2737 \$2252 \$2785 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37382 \$153 \$2808 \$1815 \$2785 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37383 \$16 \$1390 \$16 \$153 \$2785 VNB sky130_fd_sc_hd__inv_1
X$37384 \$153 \$2432 \$2377 \$2024 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37385 \$153 \$2847 \$1547 \$2884 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37386 \$16 \$1037 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37389 \$153 \$2901 \$1208 \$3037 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$37390 \$16 \$2024 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37391 \$153 \$2416 \$2377 \$1795 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37392 \$16 \$1208 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37393 \$16 \$1595 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37394 \$153 \$2885 \$1943 \$2886 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37395 \$16 \$1795 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37396 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$37397 \$16 \$1480 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37398 \$153 \$2848 \$1815 \$2886 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37400 \$153 \$2620 \$2511 \$1942 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37401 \$153 \$2849 \$2064 \$2886 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37402 \$16 \$1942 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37403 \$153 \$2850 \$1547 \$2886 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37404 \$16 \$1980 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37405 \$153 \$2809 \$2511 \$1658 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37406 \$16 \$1686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37408 \$153 \$2851 \$2887 \$1687 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37409 \$16 \$1658 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37410 \$16 \$1013 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37411 \$153 \$2810 \$2380 \$1942 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37412 \$16 \$1687 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37413 \$16 \$1404 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37414 \$16 \$1942 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37415 \$153 \$2852 \$2887 \$1658 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37417 \$153 \$2763 \$2380 \$1795 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37418 \$153 \$2852 \$1547 \$3014 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37420 \$153 \$2887 \$1553 \$2585 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$37421 \$153 \$2853 \$1815 \$3014 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37423 \$16 \$1658 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37424 \$153 \$2836 \$2646 \$1795 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37425 \$153 \$2764 \$2646 \$1658 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37426 \$153 \$2809 \$1547 \$2275 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37427 \$153 \$2739 \$1943 \$2586 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37429 \$153 \$2854 \$2064 \$2586 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37430 \$153 \$2688 \$2252 \$2586 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37431 \$153 \$2836 \$1815 \$2586 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37432 \$153 \$2764 \$1547 \$2586 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37433 \$153 \$2533 \$1792 \$1594 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37435 \$153 \$2648 \$2704 \$1942 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37436 \$16 \$1067 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37438 \$16 \$1594 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37439 \$16 \$2180 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37440 \$16 \$2006 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37441 \$153 \$2811 \$2704 \$2006 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37442 \$153 \$2633 \$2210 \$1594 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37443 \$16 \$1942 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37445 \$153 \$2811 \$1943 \$2671 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37446 \$16 \$1594 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37447 \$16 \$1795 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37448 \$16 \$1594 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37450 \$16 \$1687 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37451 \$16 \$1795 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37452 \$153 \$2812 \$2649 \$1687 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37453 \$153 \$2706 \$2649 \$1795 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37454 \$153 \$2812 \$1792 \$2741 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37456 \$16 \$2024 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37457 \$153 \$2813 \$2649 \$2024 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37460 \$153 \$2855 \$2210 \$2671 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37461 \$153 \$2814 \$2649 \$2006 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37462 \$153 \$2813 \$2210 \$2741 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37463 \$16 \$842 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37464 \$16 \$691 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37465 \$153 \$2814 \$1943 \$2741 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37466 \$16 \$2006 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37470 \$16 \$2647 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37471 \$16 \$1980 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37472 \$153 \$2689 \$1815 \$2671 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37473 \$153 \$2765 \$2649 \$1980 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37475 \$153 \$2888 \$2252 \$2889 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37476 \$153 \$2765 \$2009 \$2741 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37478 \$16 \$588 \$2647 \$2856 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$37480 \$153 \$2933 \$757 \$2856 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$37481 \$153 \$2815 \$2252 \$2743 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37482 \$153 \$2837 \$2009 \$2743 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37483 \$16 \$588 \$16 \$153 \$2889 VNB sky130_fd_sc_hd__inv_1
X$37484 \$16 \$2100 \$16 \$153 \$2674 VNB sky130_fd_sc_hd__clkbuf_2
X$37485 \$16 \$2414 \$16 \$153 \$2936 VNB sky130_fd_sc_hd__clkbuf_2
X$37486 \$153 \$2878 \$2635 \$2538 \$2674 \$2650 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$37487 \$16 \$2793 \$16 \$153 \$2100 VNB sky130_fd_sc_hd__clkbuf_2
X$37490 \$153 \$2635 \$2674 \$2816 \$2650 \$2538 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$37492 \$16 \$2729 \$16 \$153 \$1348 VNB sky130_fd_sc_hd__clkbuf_2
X$37493 \$16 \$2793 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37494 \$153 \$2857 \$1595 \$2902 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$37495 \$153 \$2674 \$2650 \$2766 \$2635 \$2538 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$37496 \$153 \$2635 \$2650 \$2786 \$2674 \$2538 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$37497 \$16 \$2816 \$16 \$153 \$1404 VNB sky130_fd_sc_hd__clkbuf_2
X$37499 \$153 \$2767 \$2652 \$2199 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37500 \$153 \$2577 \$2857 \$2199 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37501 \$153 \$2767 \$2184 \$2636 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37502 \$16 \$2199 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37503 \$153 \$2890 \$1806 \$2594 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37504 \$16 \$1965 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37507 \$16 \$2786 \$16 \$153 \$1328 VNB sky130_fd_sc_hd__clkbuf_2
X$37508 \$16 \$2199 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37509 \$16 \$945 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37510 \$16 \$1390 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37511 \$16 \$1037 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37512 \$16 \$1595 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37514 \$153 \$2744 \$2026 \$2636 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37515 \$153 \$2891 \$2026 \$2594 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37516 \$153 \$2745 \$1924 \$2636 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37517 \$16 \$757 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37519 \$153 \$2768 \$2652 \$1845 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37520 \$16 \$588 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37523 \$153 \$2678 \$2857 \$1805 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37524 \$153 \$2623 \$1703 \$2636 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37525 \$153 \$2768 \$1471 \$2636 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37526 \$153 \$2858 \$1471 \$3269 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37527 \$16 \$1845 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37528 \$16 \$1805 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37532 \$153 \$2892 \$1895 \$2879 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37533 \$153 \$2730 \$2708 \$2043 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37534 \$153 \$2893 \$1471 \$2746 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37535 \$16 \$1348 \$16 \$153 \$2746 VNB sky130_fd_sc_hd__inv_1
X$37537 \$153 \$2769 \$2708 \$1965 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37538 \$153 \$2859 \$1703 \$2879 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37540 \$16 \$2043 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37542 \$153 \$2624 \$1924 \$2746 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37543 \$153 \$2769 \$1806 \$2746 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37545 \$153 \$2838 \$2555 \$1805 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37546 \$153 \$2787 \$2184 \$2879 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37547 \$16 \$1965 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37550 \$153 \$2770 \$2555 \$1965 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37551 \$153 \$2839 \$2555 \$1923 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37552 \$153 \$2770 \$1806 \$2557 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37553 \$153 \$2838 \$1703 \$2557 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37554 \$16 \$1965 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37555 \$16 \$1923 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37556 \$153 \$2771 \$2359 \$1805 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37558 \$153 \$2860 \$2359 \$1923 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37559 \$153 \$2839 \$1895 \$2557 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37560 \$153 \$2747 \$1954 \$2327 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37561 \$16 \$2043 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37562 \$16 \$1805 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37563 \$153 \$2894 \$1471 \$2895 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37565 \$16 \$1845 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37567 \$153 \$2817 \$2525 \$1923 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37568 \$153 \$2840 \$2525 \$2089 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37569 \$16 \$1923 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37570 \$153 \$2840 \$2026 \$2499 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37571 \$16 \$2089 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37572 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$37574 \$16 \$1264 \$2347 \$2904 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$37575 \$153 \$2817 \$1895 \$2499 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37576 \$16 \$1264 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37578 \$153 \$2861 \$2597 \$2043 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37579 \$153 \$2771 \$1703 \$2327 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37580 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$37581 \$16 \$691 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37582 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$37583 \$16 \$2043 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37584 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$37586 \$153 \$2363 \$2597 \$1845 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37587 \$153 \$2862 \$2597 \$1965 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37588 \$16 \$1845 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37589 \$153 \$2862 \$1806 \$2346 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37590 \$16 \$1965 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37592 \$16 \$1805 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37593 \$153 \$2818 \$2560 \$1805 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37596 \$153 \$2880 \$2560 \$2199 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37597 \$153 \$2655 \$2560 \$2042 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37599 \$153 \$2841 \$2560 \$2043 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37602 \$16 \$2042 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37603 \$16 \$757 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37604 \$153 \$2841 \$1954 \$2637 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37605 \$153 \$2906 \$2560 \$1845 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37606 \$153 \$2749 \$1806 \$2637 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37607 \$16 \$2043 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37608 \$16 \$588 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37609 \$16 \$1845 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37610 \$16 \$588 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37611 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$37612 \$153 \$2772 \$2578 \$2199 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37614 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$37616 \$16 \$1551 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37617 \$153 \$2896 \$1703 \$2926 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37618 \$153 \$2772 \$2184 \$2500 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37619 \$16 \$1805 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37620 \$16 \$1845 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37621 \$16 \$1845 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37622 \$153 \$2714 \$2578 \$1845 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37623 \$16 \$2199 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37625 \$16 \$1965 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37627 \$153 \$2819 \$2578 \$1965 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37629 \$153 \$2819 \$1806 \$2500 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37631 \$16 \$2794 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37633 \$16 \$2820 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37634 \$16 \$2908 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37635 \$16 \$1969 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37636 \$16 \$2908 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37637 \$153 \$2122 \$2517 \$1969 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37639 \$16 \$1969 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37641 \$153 \$2864 \$2863 \$2098 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37642 \$153 \$2773 \$2517 \$2105 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37643 \$153 \$2864 \$1993 \$2639 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37645 \$153 \$2897 \$2438 \$2639 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37647 \$153 \$2821 \$2517 \$1756 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37648 \$16 \$2105 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37649 \$153 \$2863 \$1489 \$2822 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$37650 \$16 \$1044 \$1968 \$2822 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$37652 \$16 \$2016 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37653 \$16 \$1756 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37654 \$153 \$2823 \$2485 \$2016 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37656 \$16 \$2105 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37658 \$153 \$2909 \$1613 \$2639 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37659 \$16 \$1044 \$16 \$153 \$2639 VNB sky130_fd_sc_hd__inv_1
X$37661 \$153 \$2842 \$2731 \$2105 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37662 \$153 \$2751 \$1993 \$2502 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37663 \$16 \$1720 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37664 \$16 \$2774 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37665 \$16 \$1756 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37667 \$153 \$2823 \$1715 \$2502 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37668 \$153 \$2911 \$2731 \$1756 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37670 \$16 \$1878 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37671 \$153 \$2824 \$2731 \$1878 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37672 \$153 \$2842 \$2438 \$2752 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37673 \$16 \$1543 \$16 \$153 \$2752 VNB sky130_fd_sc_hd__inv_1
X$37674 \$153 \$2753 \$2731 \$2016 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37676 \$153 \$2824 \$1868 \$2752 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37677 \$153 \$2825 \$1613 \$2641 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37679 \$16 \$2104 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37680 \$153 \$2913 \$2696 \$2104 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37681 \$153 \$2788 \$1613 \$2627 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37683 \$16 \$1929 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37684 \$16 \$2232 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37685 \$16 \$1878 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37686 \$153 \$2795 \$1868 \$2627 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37687 \$153 \$2795 \$2696 \$1878 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37688 \$16 \$1760 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37689 \$16 \$1879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37690 \$153 \$2658 \$2796 \$1879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37691 \$16 \$1585 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37692 \$16 \$2659 \$16 \$153 \$2580 VNB sky130_fd_sc_hd__clkbuf_2
X$37694 \$16 \$1518 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37695 \$16 \$1811 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37696 \$16 \$2016 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37697 \$153 \$2825 \$2796 \$1969 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37698 \$153 \$2865 \$2092 \$2641 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37699 \$153 \$2683 \$2796 \$2016 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37700 \$16 \$1969 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37701 \$16 \$901 \$16 \$153 \$2641 VNB sky130_fd_sc_hd__inv_1
X$37703 \$153 \$3000 \$1868 \$2641 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37704 \$16 \$1878 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37705 \$153 \$2826 \$2866 \$1878 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37707 \$16 \$1879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37708 \$153 \$2775 \$2579 \$1879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37709 \$16 \$1879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37710 \$16 \$2462 \$2580 \$2914 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$37711 \$153 \$2826 \$1868 \$2789 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37713 \$153 \$2915 \$2866 \$1879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37714 \$153 \$2797 \$1712 \$2789 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37715 \$16 \$2462 \$16 \$153 \$2789 VNB sky130_fd_sc_hd__inv_1
X$37716 \$153 \$2775 \$1558 \$2606 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37718 \$153 \$2798 \$2881 \$1878 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37721 \$16 \$2462 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37723 \$16 \$1756 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37724 \$153 \$2798 \$1868 \$2790 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37725 \$153 \$2867 \$2881 \$1969 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37726 \$153 \$2799 \$1558 \$2790 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37727 \$16 \$1184 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37728 \$16 \$1969 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37731 \$153 \$2881 \$700 \$2800 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$37733 \$153 \$2867 \$1613 \$2790 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37734 \$16 \$815 \$16 \$153 \$2790 VNB sky130_fd_sc_hd__inv_1
X$37736 \$16 \$815 \$2580 \$2800 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$37737 \$153 \$2868 \$2916 \$1969 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37738 \$16 \$1969 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37739 \$16 \$2580 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37740 \$16 \$700 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37741 \$16 \$815 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37744 \$16 \$2016 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37745 \$153 \$2843 \$2732 \$1879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37746 \$153 \$2801 \$2092 \$2791 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37747 \$153 \$2776 \$2732 \$2016 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37748 \$153 \$2882 \$1993 \$2791 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37749 \$16 \$2580 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37750 \$153 \$2777 \$2732 \$1756 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37752 \$16 \$1120 \$2580 \$2869 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$37753 \$153 \$2916 \$1303 \$2869 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$37754 \$153 \$2777 \$1712 \$2504 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37755 \$16 \$1120 \$16 \$153 \$2791 VNB sky130_fd_sc_hd__inv_1
X$37756 \$16 \$2827 \$16 \$153 \$1543 VNB sky130_fd_sc_hd__clkbuf_2
X$37757 \$16 \$2189 \$16 \$153 \$2685 VNB sky130_fd_sc_hd__clkbuf_2
X$37758 \$153 \$2917 \$2699 \$2733 \$2684 \$2685 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$37760 \$153 \$2827 \$2684 \$2733 \$2699 \$2685 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$37761 \$16 \$2733 \$2685 \$2699 \$2684 \$16 \$153 \$2898 VNB
+ sky130_fd_sc_hd__and4_2
X$37762 \$16 \$1303 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37764 \$153 \$2754 \$2684 \$2699 \$2685 \$2733 \$16 \$16 VNB
+ sky130_fd_sc_hd__nor4b_2
X$37765 \$153 \$2684 \$2685 \$2792 \$2699 \$2733 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$37766 \$16 \$1044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37768 \$16 \$1489 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37769 \$153 \$2802 \$1936 \$2613 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37771 \$16 \$1972 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37772 \$153 \$2828 \$2271 \$2613 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37773 \$153 \$2828 \$2612 \$2085 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37774 \$153 \$2870 \$2267 \$2899 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37776 \$153 \$2802 \$2612 \$2031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37777 \$16 \$2792 \$16 \$153 \$1475 VNB sky130_fd_sc_hd__clkbuf_2
X$37779 \$153 \$2829 \$1936 \$2899 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37780 \$16 \$2031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37781 \$16 \$2898 \$16 \$153 \$1585 VNB sky130_fd_sc_hd__clkbuf_2
X$37782 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$37783 \$16 \$2191 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37784 \$153 \$2871 \$2056 \$2899 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37785 \$153 \$2778 \$2612 \$2192 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37787 \$16 \$1585 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37790 \$16 \$2192 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37791 \$153 \$2830 \$2612 \$1860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37792 \$153 \$2702 \$2086 \$2613 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37793 \$16 \$1960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37794 \$16 \$1860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37795 \$16 \$2093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37796 \$153 \$2918 \$2831 \$2093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37797 \$153 \$2778 \$2269 \$2613 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37799 \$153 \$2831 \$1245 \$2756 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$37800 \$16 \$2232 \$16 \$153 \$2872 VNB sky130_fd_sc_hd__inv_1
X$37802 \$16 \$1960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37803 \$153 \$2919 \$2831 \$1960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37804 \$153 \$2832 \$998 \$2779 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$37805 \$16 \$998 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37808 \$16 \$2031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37809 \$16 \$2803 \$16 \$153 \$1972 VNB sky130_fd_sc_hd__clkbuf_2
X$37810 \$16 \$901 \$16 \$153 \$2780 VNB sky130_fd_sc_hd__inv_1
X$37811 \$153 \$2873 \$2832 \$1860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37812 \$153 \$2833 \$2581 \$2031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37813 \$153 \$2833 \$1936 \$2491 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37814 \$16 \$2803 \$16 \$153 \$1885 VNB sky130_fd_sc_hd__clkbuf_2
X$37817 \$16 \$2031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37818 \$16 \$2803 \$16 \$153 \$2531 VNB sky130_fd_sc_hd__clkbuf_2
X$37820 \$16 \$2085 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37821 \$153 \$2781 \$2581 \$2085 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37822 \$16 \$1973 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37823 \$153 \$2834 \$2832 \$1973 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37824 \$153 \$2758 \$2267 \$2491 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37825 \$16 \$2462 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37826 \$16 \$2093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37829 \$16 \$2462 \$16 \$153 \$2920 VNB sky130_fd_sc_hd__inv_1
X$37830 \$16 \$2192 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37831 \$153 \$2662 \$2570 \$2192 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37832 \$153 \$2875 \$2874 \$2093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37833 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$37834 \$153 \$2875 \$2265 \$2920 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37836 \$16 \$2093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37838 \$153 \$2782 \$2570 \$2093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37839 \$153 \$2876 \$2570 \$2085 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37840 \$153 \$2876 \$2271 \$2508 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37841 \$153 \$2782 \$2265 \$2508 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37844 \$16 \$815 \$2531 \$2783 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$37846 \$16 \$700 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37847 \$16 \$2192 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37848 \$153 \$2760 \$2804 \$2192 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37850 \$16 \$1973 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37851 \$153 \$2922 \$2804 \$1973 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37852 \$16 \$1860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37853 \$16 \$1120 \$2531 \$2784 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$37855 \$153 \$2761 \$2804 \$2031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37857 \$153 \$2835 \$2804 \$1860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37858 \$16 \$2031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37859 \$153 \$2883 \$1303 \$2784 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$37860 \$153 \$2835 \$2000 \$2759 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37861 \$16 \$2093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37864 \$153 \$2762 \$2572 \$2085 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37865 \$16 \$2085 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37866 \$153 \$2495 \$2271 \$2032 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37867 \$153 \$2900 \$2265 \$2642 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37869 \$16 \$1860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37870 \$153 \$2805 \$2271 \$2642 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37871 \$153 \$2877 \$2883 \$2191 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37873 \$153 \$2509 \$2572 \$1860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37875 \$16 \$1973 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37876 \$153 \$2667 \$2883 \$1973 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37878 \$153 \$2806 \$2000 \$2642 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37879 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$37884 \$16 \$1960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37885 \$16 \$2192 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37886 \$153 \$2844 \$2883 \$1960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37887 \$153 \$2617 \$2572 \$2192 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37888 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$37890 \$153 \$3055 \$1936 \$2923 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37893 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$37894 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$37895 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$37896 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$37897 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$37898 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$37899 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$37900 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$37901 \$153 \$6139 \$6178 \$5181 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37903 \$153 \$6219 \$6178 \$5245 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37905 \$153 \$6139 \$5174 \$6174 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37906 \$16 \$5245 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37909 \$153 \$6219 \$5107 \$6174 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37911 \$16 \$4742 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37912 \$16 \$4742 \$6051 \$6207 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$37914 \$153 \$6178 \$5152 \$6207 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$37915 \$153 \$6140 \$6178 \$5274 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37916 \$16 \$5152 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37917 \$16 \$5274 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37919 \$153 \$6140 \$4706 \$6174 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37920 \$153 \$6220 \$6178 \$5404 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37921 \$153 \$5536 \$5373 \$4579 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37922 \$153 \$6220 \$5177 \$6174 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37923 \$16 \$4742 \$16 \$153 \$6174 VNB sky130_fd_sc_hd__inv_1
X$37924 \$16 \$5489 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37925 \$16 \$5403 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37926 \$153 \$6141 \$5976 \$5403 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37927 \$16 \$5404 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37929 \$153 \$5992 \$5976 \$5736 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37930 \$153 \$6141 \$5405 \$5977 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37931 \$153 \$6258 \$5405 \$6257 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37932 \$16 \$5080 \$6051 \$6276 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$37933 \$16 \$5736 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37936 \$153 \$6277 \$6251 \$5274 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37937 \$16 \$5181 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37938 \$16 \$5274 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37939 \$153 \$6052 \$5976 \$5404 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37940 \$153 \$6259 \$5107 \$6260 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37941 \$16 \$5404 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37942 \$16 \$5181 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37943 \$16 \$5080 \$16 \$153 \$6260 VNB sky130_fd_sc_hd__inv_1
X$37944 \$153 \$6126 \$6053 \$5181 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37947 \$153 \$6054 \$6053 \$5489 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37948 \$153 \$6208 \$6053 \$5518 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37949 \$153 \$6179 \$6053 \$5404 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37951 \$16 \$5518 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37952 \$153 \$6179 \$5177 \$6043 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37953 \$16 \$4896 \$6051 \$6278 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$37955 \$153 \$6127 \$6056 \$5518 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37956 \$153 \$6209 \$6056 \$5245 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37957 \$16 \$5518 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37958 \$16 \$5245 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37960 \$16 \$6051 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37961 \$16 \$4812 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37962 \$16 \$6051 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37963 \$153 \$6142 \$6056 \$5489 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37964 \$16 \$5736 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37965 \$153 \$6128 \$6056 \$5736 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37966 \$153 \$6142 \$5373 \$5993 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37967 \$16 \$4947 \$6051 \$6279 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$37968 \$16 \$5181 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37970 \$153 \$5947 \$5405 \$5993 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37971 \$153 \$6221 \$5948 \$5181 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37972 \$16 \$5489 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37973 \$16 \$4947 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37975 \$153 \$6180 \$5373 \$6143 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37976 \$153 \$6221 \$5174 \$6143 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37977 \$16 \$5274 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37979 \$16 \$5026 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37980 \$16 \$4600 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37982 \$153 \$6182 \$5948 \$5736 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37983 \$153 \$6181 \$5463 \$6143 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37984 \$153 \$6144 \$5107 \$6143 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37986 \$153 \$6281 \$5874 \$5404 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37987 \$153 \$6182 \$5055 \$6143 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37989 \$153 \$6129 \$5874 \$5181 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37991 \$153 \$6222 \$5874 \$5518 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37992 \$153 \$6210 \$5874 \$5736 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$37993 \$16 \$5404 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37994 \$16 \$5518 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37995 \$16 \$5026 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$37997 \$153 \$6210 \$5055 \$5890 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37998 \$153 \$6222 \$5463 \$5890 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$37999 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$38000 \$16 \$5736 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38002 \$16 \$5736 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38004 \$153 \$6261 \$5107 \$6044 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38005 \$153 \$6145 \$5055 \$6044 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38006 \$16 \$5181 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38010 \$153 \$6211 \$6120 \$5404 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38011 \$16 \$4712 \$5630 \$6223 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$38013 \$153 \$6211 \$5177 \$6044 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38014 \$153 \$6224 \$5373 \$6044 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38015 \$16 \$5404 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38017 \$153 \$6130 \$6060 \$5274 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38018 \$16 \$4712 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38019 \$16 \$5404 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38021 \$153 \$6283 \$6060 \$5404 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38022 \$153 \$6183 \$5373 \$6045 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38023 \$16 \$5181 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38025 \$153 \$6284 \$6060 \$5181 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38027 \$153 \$6184 \$5055 \$6177 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38030 \$153 \$6146 \$5405 \$6045 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38031 \$153 \$6285 \$6060 \$5736 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38032 \$16 \$4742 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38033 \$16 \$5152 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38034 \$153 \$6121 \$5152 \$6185 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$38035 \$16 \$4742 \$5900 \$6185 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$38036 \$16 \$5736 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38037 \$16 \$5900 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38039 \$153 \$6225 \$6121 \$5271 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38040 \$153 \$6148 \$6121 \$5324 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38043 \$153 \$6225 \$5069 \$6149 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38044 \$153 \$6147 \$5406 \$6149 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38045 \$153 \$6226 \$6121 \$5478 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38047 \$153 \$6148 \$5096 \$6149 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38048 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$38049 \$153 \$6226 \$5390 \$6149 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38050 \$153 \$6186 \$6121 \$5232 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38051 \$16 \$5478 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38052 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$38054 \$16 \$5051 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38055 \$16 \$5232 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38056 \$153 \$6131 \$6121 \$5469 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38057 \$153 \$6186 \$5205 \$6149 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38058 \$153 \$6287 \$5051 \$6187 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$38059 \$16 \$5080 \$5900 \$6187 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$38060 \$16 \$5469 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38062 \$153 \$6227 \$6287 \$5271 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38063 \$16 \$5900 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38064 \$153 \$6189 \$6287 \$5338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38066 \$153 \$6227 \$5069 \$6262 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38067 \$153 \$6188 \$5096 \$6262 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38068 \$16 \$5271 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38070 \$16 \$5338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38072 \$16 \$5080 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38074 \$153 \$6190 \$5846 \$5478 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38075 \$153 \$6150 \$5846 \$5232 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38077 \$16 \$5232 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38078 \$153 \$6150 \$5205 \$6032 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38079 \$16 \$5478 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38080 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$38081 \$153 \$6263 \$5209 \$6264 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38083 \$153 \$6190 \$5390 \$6032 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38084 \$153 \$6191 \$5846 \$5469 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38085 \$153 \$6062 \$5096 \$6032 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38087 \$153 \$6191 \$5287 \$6032 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38088 \$16 \$5469 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38090 \$16 \$4947 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38094 \$153 \$6151 \$5849 \$5232 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38095 \$153 \$6132 \$5849 \$5478 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38096 \$153 \$6151 \$5205 \$5980 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38097 \$16 \$5232 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38098 \$16 \$5478 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38099 \$16 \$5900 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38101 \$153 \$6289 \$5849 \$5566 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38104 \$153 \$6192 \$5849 \$5469 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38105 \$153 \$6194 \$5929 \$5566 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38106 \$153 \$6192 \$5287 \$5980 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38107 \$16 \$5469 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38108 \$16 \$5566 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38110 \$153 \$6228 \$5929 \$5478 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38111 \$16 \$5338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38112 \$153 \$6193 \$5929 \$5338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38113 \$153 \$6228 \$5390 \$5852 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38114 \$153 \$6193 \$5209 \$5852 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38115 \$153 \$6229 \$6001 \$5338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38117 \$153 \$6194 \$5519 \$5852 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38118 \$16 \$5026 \$5479 \$6152 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$38119 \$153 \$6229 \$5209 \$6122 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38120 \$16 \$4600 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38122 \$153 \$6212 \$6123 \$5232 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38123 \$16 \$5338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38124 \$16 \$5026 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38125 \$16 \$4822 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38128 \$16 \$4494 \$16 \$153 \$6291 VNB sky130_fd_sc_hd__inv_1
X$38129 \$153 \$6133 \$6123 \$5469 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38130 \$153 \$6212 \$5205 \$5982 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38131 \$16 \$4822 \$5479 \$6292 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$38132 \$16 \$5271 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38133 \$153 \$6134 \$6123 \$5566 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38134 \$16 \$5232 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38135 \$16 \$5271 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38136 \$16 \$5469 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38139 \$153 \$6213 \$6123 \$5338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38140 \$153 \$6213 \$5209 \$5982 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38141 \$16 \$5338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38142 \$16 \$5566 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38143 \$153 \$6153 \$6085 \$5478 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38144 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$38146 \$16 \$5566 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38148 \$153 \$6294 \$6085 \$5566 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38150 \$153 \$6153 \$5390 \$6175 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38151 \$153 \$6154 \$5406 \$6175 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38152 \$16 \$4869 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38154 \$16 \$5271 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38155 \$153 \$6230 \$6085 \$5271 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38156 \$16 \$5478 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38159 \$153 \$6155 \$6085 \$5469 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38160 \$153 \$6230 \$5069 \$6175 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38161 \$153 \$6155 \$5287 \$6175 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38163 \$153 \$6231 \$6200 \$6136 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38164 \$153 \$6214 \$6195 \$5605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38166 \$153 \$6231 \$6195 \$5819 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38167 \$153 \$6156 \$5775 \$6005 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38168 \$153 \$6069 \$6195 \$5702 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38169 \$16 \$5796 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38170 \$16 \$5605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38171 \$16 \$5714 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38173 \$153 \$6086 \$5755 \$6005 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38175 \$153 \$6197 \$6195 \$5834 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38176 \$153 \$6196 \$5775 \$6136 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38177 \$16 \$4760 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38178 \$153 \$6197 \$5881 \$6136 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38179 \$16 \$5834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38181 \$16 \$4760 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38182 \$16 \$5452 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38184 \$16 \$5528 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38185 \$153 \$6265 \$5452 \$6297 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$38186 \$153 \$6157 \$6195 \$5528 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38187 \$16 \$4780 \$5428 \$6232 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$38188 \$153 \$6157 \$5500 \$6136 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38190 \$153 \$6266 \$5795 \$6267 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38192 \$16 \$5528 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38194 \$16 \$4930 \$16 \$153 \$6267 VNB sky130_fd_sc_hd__inv_1
X$38195 \$153 \$6158 \$5961 \$5528 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38196 \$153 \$6198 \$5961 \$5605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38198 \$153 \$6158 \$5500 \$5891 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38199 \$16 \$5605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38200 \$16 \$5259 \$6252 \$6233 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$38202 \$153 \$6198 \$5625 \$5891 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38204 \$153 \$6333 \$5543 \$6233 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$38205 \$16 \$5259 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38206 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$38207 \$16 \$5259 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38208 \$16 \$5543 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38209 \$153 \$6268 \$5755 \$6234 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38211 \$153 \$6159 \$5755 \$5891 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38212 \$16 \$5259 \$16 \$153 \$6234 VNB sky130_fd_sc_hd__inv_1
X$38214 \$16 \$1433 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38215 \$16 \$1433 \$16 \$153 \$6124 VNB sky130_fd_sc_hd__clkbuf_2
X$38217 \$16 \$5819 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38218 \$153 \$6160 \$5973 \$5819 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38219 \$16 \$5819 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38220 \$16 \$5834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38221 \$153 \$6199 \$5973 \$5834 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38222 \$153 \$6160 \$6200 \$6089 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38223 \$16 \$6124 \$16 \$153 \$6252 VNB sky130_fd_sc_hd__clkbuf_2
X$38225 \$153 \$6199 \$5881 \$6089 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38226 \$153 \$6235 \$6253 \$5702 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38228 \$153 \$6161 \$5973 \$5856 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38229 \$16 \$5856 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38230 \$16 \$5702 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38232 \$16 \$5834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38233 \$153 \$6236 \$6253 \$5834 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38236 \$153 \$6161 \$5795 \$6089 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38237 \$16 \$5819 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38238 \$16 \$5796 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38239 \$153 \$6235 \$5470 \$6421 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38240 \$153 \$6163 \$6011 \$5796 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38241 \$16 \$4562 \$16 \$153 \$6421 VNB sky130_fd_sc_hd__inv_1
X$38242 \$16 \$4882 \$6269 \$6237 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$38244 \$153 \$6238 \$4781 \$6237 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$38245 \$153 \$6162 \$6200 \$5985 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38246 \$153 \$6163 \$5775 \$5985 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38247 \$16 \$5834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38248 \$16 \$6269 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38249 \$16 \$4781 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38250 \$16 \$6124 \$16 \$153 \$5906 VNB sky130_fd_sc_hd__clkbuf_2
X$38252 \$16 \$5819 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38253 \$16 \$5528 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38254 \$153 \$6270 \$5795 \$6176 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38255 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$38257 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$38258 \$153 \$6164 \$5470 \$5985 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38260 \$153 \$6239 \$6238 \$5819 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38261 \$153 \$6201 \$5755 \$6176 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38262 \$16 \$4882 \$16 \$153 \$6176 VNB sky130_fd_sc_hd__inv_1
X$38263 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$38264 \$16 \$4882 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38265 \$16 \$5819 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38268 \$153 \$6300 \$5500 \$5892 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38269 \$153 \$6202 \$6012 \$5819 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38270 \$153 \$6202 \$6200 \$5892 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38271 \$153 \$6203 \$6012 \$5856 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38273 \$153 \$6203 \$5795 \$5892 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38276 \$153 \$6070 \$5775 \$5892 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38277 \$16 \$5856 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38278 \$16 \$5799 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38279 \$16 \$5834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38280 \$16 \$5400 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38281 \$16 \$5819 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38283 \$153 \$6240 \$6271 \$5819 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38284 \$16 \$5819 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38285 \$153 \$6165 \$6072 \$5819 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38287 \$153 \$6241 \$6271 \$5856 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38289 \$153 \$6165 \$6200 \$5987 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38290 \$153 \$6271 \$4784 \$6204 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$38291 \$153 \$6242 \$6271 \$5605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38293 \$16 \$4567 \$5906 \$6204 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$38294 \$16 \$5605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38295 \$153 \$6166 \$6072 \$5714 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38297 \$153 \$6243 \$6271 \$5714 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38298 \$153 \$6166 \$5755 \$5987 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38299 \$16 \$4567 \$16 \$153 \$6318 VNB sky130_fd_sc_hd__inv_1
X$38300 \$16 \$4567 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38302 \$153 \$6243 \$5755 \$6318 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38303 \$16 \$4567 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38305 \$153 \$6075 \$5907 \$5887 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38306 \$16 \$4930 \$6216 \$6272 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$38307 \$16 \$4930 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38308 \$153 \$6254 \$5484 \$6273 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38309 \$16 \$5887 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38311 \$16 \$5452 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38312 \$16 \$4590 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38313 \$153 \$6244 \$5452 \$6303 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$38316 \$16 \$4780 \$5485 \$6205 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$38317 \$153 \$6076 \$4590 \$6205 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$38318 \$153 \$6074 \$5938 \$5823 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38319 \$16 \$5786 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38320 \$16 \$5636 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38321 \$16 \$4760 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38322 \$153 \$6215 \$6076 \$5636 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38323 \$16 \$5609 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38324 \$16 \$5963 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38326 \$153 \$6137 \$6076 \$5963 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38327 \$16 \$5786 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38328 \$153 \$6046 \$6076 \$5609 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38329 \$153 \$6245 \$6076 \$5786 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38331 \$153 \$6167 \$6076 \$5887 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38332 \$153 \$6245 \$5635 \$6018 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38333 \$153 \$6206 \$5543 \$6305 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$38334 \$153 \$6167 \$5627 \$6018 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38335 \$153 \$6168 \$6206 \$5579 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38338 \$153 \$6079 \$6206 \$5786 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38339 \$153 \$6168 \$5484 \$6047 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38340 \$153 \$6246 \$6206 \$5887 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38341 \$16 \$6078 \$16 \$153 \$6216 VNB sky130_fd_sc_hd__clkbuf_2
X$38342 \$16 \$5579 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38344 \$153 \$6080 \$6169 \$5786 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38345 \$153 \$6246 \$5627 \$6047 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38346 \$16 \$5259 \$16 \$153 \$6047 VNB sky130_fd_sc_hd__inv_1
X$38347 \$16 \$5786 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38348 \$16 \$5963 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38350 \$16 \$5259 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38351 \$153 \$6306 \$5806 \$6048 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38352 \$16 \$5636 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38353 \$153 \$6138 \$6169 \$5636 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38355 \$153 \$6247 \$6169 \$5718 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38356 \$16 \$5786 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38357 \$153 \$6170 \$5835 \$5786 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38358 \$16 \$5718 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38359 \$16 \$4882 \$6255 \$6248 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$38360 \$153 \$6308 \$4781 \$6248 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$38362 \$16 \$5963 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38363 \$153 \$6170 \$5635 \$5867 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38364 \$153 \$6247 \$5938 \$6048 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38366 \$153 \$6217 \$5910 \$5718 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38367 \$153 \$6081 \$5074 \$6048 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38370 \$16 \$5767 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38371 \$153 \$6217 \$5938 \$5893 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38372 \$153 \$6171 \$5910 \$5767 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38373 \$153 \$6249 \$5910 \$5786 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38374 \$153 \$6171 \$5575 \$5893 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38375 \$153 \$6249 \$5635 \$5893 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38379 \$16 \$5963 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38380 \$153 \$6082 \$5941 \$5963 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38381 \$153 \$6310 \$5627 \$5893 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38382 \$153 \$6312 \$5938 \$6311 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38383 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$38386 \$16 \$5609 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38387 \$16 \$4963 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38388 \$153 \$6172 \$5941 \$5609 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38391 \$16 \$4784 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38392 \$153 \$5012 \$3893 \$4963 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38393 \$153 \$6256 \$4784 \$6313 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$38394 \$153 \$6172 \$5074 \$5894 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38395 \$16 \$4376 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38397 \$16 \$5718 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38400 \$153 \$6250 \$5938 \$6274 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38401 \$16 \$5767 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38402 \$153 \$6173 \$6023 \$5767 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38403 \$153 \$6250 \$6256 \$5718 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38404 \$153 \$6173 \$5575 \$5895 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38405 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$38406 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$38408 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$38409 \$16 \$5636 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38410 \$16 \$5609 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38411 \$153 \$6314 \$6023 \$5609 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38412 \$153 \$6218 \$6023 \$5636 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38413 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$38414 \$153 \$6218 \$5509 \$5895 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38416 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$38417 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$38418 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$38419 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$38420 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$38421 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$38422 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$38423 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$38424 \$153 \$3588 \$3494 \$3766 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38425 \$153 \$3472 \$3494 \$3474 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38426 \$16 \$3474 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38427 \$16 \$3766 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38428 \$153 \$3472 \$3490 \$3420 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38429 \$16 \$3709 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38432 \$153 \$3550 \$3494 \$3385 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38433 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$38434 \$153 \$3513 \$3494 \$3473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38435 \$16 \$3385 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38436 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$38438 \$153 \$3513 \$3540 \$3420 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38439 \$16 \$3473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38442 \$153 \$3421 \$3494 \$3571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38443 \$16 \$3615 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38445 \$16 \$3692 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38446 \$16 \$3686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38448 \$153 \$3330 \$3495 \$3385 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38449 \$153 \$3514 \$3495 \$3474 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38451 \$16 \$3385 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38452 \$153 \$3514 \$3490 \$3331 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38453 \$153 \$3423 \$3495 \$3473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38455 \$153 \$3496 \$3495 \$3571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38456 \$16 \$3474 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38457 \$16 \$3473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38458 \$16 \$2024 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38461 \$16 \$3571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38462 \$153 \$3496 \$3422 \$3331 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38463 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$38464 \$153 \$3425 \$3497 \$3571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38465 \$153 \$3515 \$3497 \$3473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38466 \$16 \$3571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38468 \$153 \$3498 \$3497 \$3474 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38471 \$153 \$3515 \$3540 \$3426 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38472 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$38473 \$153 \$3498 \$3490 \$3426 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38475 \$153 \$3577 \$3407 \$3473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38476 \$16 \$3474 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38477 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$38479 \$153 \$3427 \$3407 \$3385 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38480 \$153 \$3577 \$3540 \$3578 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38481 \$16 \$3473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38483 \$16 \$3385 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38484 \$153 \$3428 \$3407 \$3474 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38486 \$153 \$3579 \$3478 \$3578 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38488 \$16 \$3766 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38489 \$16 \$3714 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38490 \$16 \$3474 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38491 \$16 \$3686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38492 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$38494 \$153 \$3475 \$3408 \$3474 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38495 \$153 \$3551 \$3408 \$3473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38496 \$16 \$3474 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38497 \$16 \$3473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38499 \$153 \$3429 \$3408 \$3385 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38501 \$153 \$3475 \$3490 \$3476 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38502 \$153 \$3447 \$3422 \$3476 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38503 \$153 \$3551 \$3540 \$3476 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38505 \$153 \$3430 \$3499 \$3473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38506 \$16 \$3385 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38507 \$16 \$3615 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38510 \$153 \$3552 \$3499 \$3571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38511 \$16 \$3473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38512 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$38513 \$153 \$3477 \$3499 \$3474 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38514 \$153 \$3552 \$3422 \$3409 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38515 \$16 \$3571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38516 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$38518 \$153 \$3477 \$3490 \$3409 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38519 \$153 \$3395 \$3410 \$3474 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38521 \$16 \$3491 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38522 \$153 \$3491 \$2024 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$38523 \$16 \$3474 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38524 \$16 \$1551 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38525 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$38527 \$153 \$3590 \$3410 \$3473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38528 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$38529 \$153 \$1407 \$3385 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$38530 \$16 \$3473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38531 \$153 \$1625 \$3473 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$38533 \$16 \$1407 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38535 \$153 \$1775 \$3474 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$38536 \$153 \$3580 \$3422 \$3334 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38537 \$153 \$3304 \$2210 \$2743 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38538 \$16 \$1775 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38540 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38542 \$153 \$1610 \$3766 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$38543 \$153 \$1538 \$3615 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$38544 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38545 \$153 \$3553 \$1482 \$1943 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38546 \$16 \$3384 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38547 \$16 \$3384 \$16 \$153 \$2233 VNB sky130_fd_sc_hd__clkbuf_2
X$38549 \$153 \$3040 \$2252 \$2634 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38550 \$153 \$3095 \$2009 \$2634 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38552 \$153 \$3479 \$1482 \$3389 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38553 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38554 \$16 \$1610 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38556 \$16 \$3389 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38557 \$153 \$3591 \$3541 \$3237 \$3554 \$3555 \$3411 \$3592 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$38559 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38560 \$153 \$3414 \$1482 \$3606 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38561 \$16 \$3606 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38562 \$153 \$3581 \$3412 \$3572 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38563 \$16 \$2634 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38564 \$16 \$3516 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38567 \$16 \$3411 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38569 \$153 \$3451 \$3079 \$3336 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38570 \$153 \$3581 \$3101 \$3336 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38571 \$153 \$3500 \$3412 \$3480 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38572 \$153 \$3582 \$3556 \$3336 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38575 \$153 \$3500 \$3504 \$3336 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38576 \$153 \$3432 \$3412 \$3386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38578 \$153 \$3517 \$3713 \$3480 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38579 \$16 \$3480 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38580 \$16 \$3386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38581 \$16 \$3687 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38582 \$153 \$3517 \$3504 \$3583 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38583 \$16 \$3480 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38585 \$153 \$3518 \$3713 \$3386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38586 \$153 \$3501 \$3713 \$3492 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38587 \$153 \$3501 \$3354 \$3583 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38588 \$153 \$3518 \$3435 \$3583 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38589 \$153 \$3348 \$3502 \$3492 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38591 \$153 \$3503 \$3502 \$3480 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38592 \$153 \$3503 \$3504 \$3337 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38593 \$153 \$3338 \$3502 \$3573 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38594 \$16 \$3480 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38595 \$16 \$3492 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38598 \$153 \$3350 \$3413 \$3492 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38599 \$16 \$3573 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38600 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$38601 \$153 \$3505 \$3413 \$3573 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38602 \$16 \$3492 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38603 \$153 \$3519 \$3413 \$3480 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38606 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38607 \$153 \$3519 \$3504 \$3339 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38608 \$16 \$3480 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38609 \$16 \$3573 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38610 \$16 \$3478 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38611 \$153 \$3520 \$3542 \$3492 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38612 \$153 \$3557 \$1482 \$3478 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38615 \$153 \$3505 \$3079 \$3339 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38616 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38617 \$153 \$3520 \$3354 \$3506 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38619 \$153 \$3481 \$1482 \$3307 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38620 \$153 \$3558 \$3542 \$3386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38621 \$153 \$3521 \$3542 \$3573 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38624 \$153 \$3558 \$3435 \$3506 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38625 \$16 \$3543 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38626 \$16 \$3386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38627 \$153 \$3521 \$3079 \$3506 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38629 \$153 \$3433 \$3493 \$3573 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38630 \$16 \$3573 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38631 \$16 \$1294 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38634 \$16 \$1597 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38635 \$153 \$3434 \$3493 \$3386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38637 \$153 \$3353 \$3493 \$3492 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38638 \$16 \$3386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38639 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$38640 \$16 \$3492 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38641 \$16 \$3573 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38642 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$38643 \$153 \$3482 \$3574 \$3480 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38645 \$153 \$3507 \$3574 \$3572 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38646 \$153 \$3507 \$3101 \$3436 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38647 \$153 \$3437 \$3574 \$3492 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38648 \$16 \$3572 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38649 \$16 \$3480 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38653 \$16 \$3386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38655 \$16 \$3509 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38656 \$153 \$3453 \$3435 \$3436 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38657 \$153 \$3508 \$2043 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$38658 \$16 \$3492 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38659 \$16 \$3344 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38660 \$16 \$3508 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38661 \$153 \$3584 \$3435 \$3585 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38662 \$153 \$3812 \$3354 \$3585 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38665 \$153 \$3373 \$2042 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$38666 \$153 \$153 \$1954 \$3292 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38667 \$153 \$153 \$2184 \$3292 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38668 \$153 \$3559 \$1482 \$1895 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38669 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38672 \$153 \$153 \$1471 \$3292 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38673 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38674 \$153 \$3356 \$1482 \$3608 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38675 \$153 \$3456 \$1482 \$1954 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38676 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38678 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38680 \$153 \$3560 \$1482 \$1471 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38682 \$153 \$3491 \$2105 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$38683 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38684 \$153 \$3770 \$1482 \$2092 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38685 \$16 \$3491 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38686 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38687 \$16 \$3241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38689 \$16 \$3272 \$3509 \$3202 \$695 \$16 \$153 VNB sky130_fd_sc_hd__mux2_1
X$38690 \$153 \$3618 \$1482 \$1993 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38691 \$153 \$3288 \$1756 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$38692 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38693 \$16 \$3288 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38694 \$16 \$3556 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38696 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38697 \$153 \$3483 \$1482 \$2026 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38699 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38701 \$153 \$3522 \$3281 \$1878 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38702 \$16 \$3310 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38703 \$153 \$3544 \$2438 \$3341 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38704 \$153 \$3544 \$3281 \$2105 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38706 \$153 \$3522 \$1868 \$3341 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38708 \$153 \$3595 \$3281 \$2016 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38709 \$16 \$2104 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38710 \$153 \$3523 \$3281 \$2104 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38711 \$16 \$2016 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38712 \$16 \$3418 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38714 \$153 \$3523 \$2092 \$3341 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38716 \$16 \$2104 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38717 \$153 \$3524 \$3211 \$1756 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38719 \$16 \$1878 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38720 \$153 \$3561 \$3211 \$1878 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38721 \$16 \$1756 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38722 \$16 \$2935 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38723 \$16 \$1543 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38726 \$153 \$3375 \$1993 \$3203 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38727 \$16 \$1628 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38728 \$16 \$1566 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38730 \$16 \$1878 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38731 \$153 \$3484 \$3282 \$1878 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38732 \$153 \$3561 \$1868 \$3203 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38733 \$153 \$3524 \$1712 \$3203 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38734 \$153 \$3485 \$3282 \$2105 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38737 \$153 \$3596 \$3282 \$2016 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38738 \$153 \$3485 \$2438 \$3246 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38739 \$16 \$2105 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38740 \$153 \$3545 \$3140 \$2105 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38741 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$38742 \$16 \$1878 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38744 \$153 \$3486 \$3140 \$1878 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38745 \$153 \$3562 \$3140 \$1756 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38746 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$38747 \$16 \$2105 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38748 \$153 \$3525 \$3225 \$2105 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38749 \$16 \$1756 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38750 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$38752 \$16 \$2016 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38753 \$153 \$3405 \$1712 \$3317 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38754 \$16 \$1878 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38755 \$153 \$3563 \$3225 \$2016 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38756 \$153 \$3526 \$3225 \$1878 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38757 \$16 \$3731 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38759 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$38760 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$38761 \$16 \$2104 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38762 \$16 \$2016 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38763 \$153 \$3487 \$3283 \$2104 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38764 \$153 \$3438 \$3283 \$2016 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38765 \$153 \$3487 \$2092 \$3131 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38766 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$38767 \$16 \$2105 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38769 \$16 \$1878 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38771 \$153 \$3488 \$3283 \$1878 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38772 \$153 \$3564 \$3283 \$2105 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38773 \$153 \$3488 \$1868 \$3131 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38774 \$153 \$3564 \$2438 \$3131 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38776 \$153 \$3527 \$3322 \$1969 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38777 \$16 \$1969 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38779 \$16 \$3560 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38780 \$16 \$4049 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38781 \$153 \$3530 \$3528 \$3560 \$4049 \$3575 \$3532 \$3511 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$38782 \$153 \$3458 \$2092 \$3296 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38784 \$153 \$3530 \$3529 \$3483 \$4223 \$3510 \$3377 \$3511 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$38786 \$153 \$3527 \$1613 \$3296 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38787 \$16 \$3598 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38788 \$16 \$3599 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38790 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38791 \$153 \$3547 \$1482 \$3565 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38792 \$153 \$3376 \$1712 \$3296 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38794 \$153 \$3530 \$3088 \$3402 \$4408 \$3547 \$3459 \$3511 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$38795 \$153 \$3530 \$3184 \$3546 \$3576 \$3548 \$3531 \$3511 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$38797 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38798 \$153 \$3532 \$1482 \$1936 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38799 \$16 \$3546 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38802 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38803 \$153 \$3548 \$1482 \$3142 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38804 \$153 \$3531 \$1482 \$2269 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38805 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38807 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38808 \$153 \$3566 \$1482 \$2086 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38810 \$153 \$3533 \$1482 \$2271 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38811 \$16 \$2086 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38812 \$16 \$3142 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38813 \$16 \$3508 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38814 \$16 \$2271 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38815 \$16 \$2265 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38816 \$16 \$3719 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38817 \$153 \$3927 \$4414 \$3586 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38819 \$153 \$3460 \$2265 \$3186 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38821 \$153 \$3378 \$2271 \$3186 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38822 \$16 \$3461 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38823 \$16 \$3461 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38824 \$153 \$3363 \$3185 \$1860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38825 \$16 \$3461 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38826 \$16 \$3461 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38827 \$16 \$3567 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38828 \$16 \$3602 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38829 \$153 \$3587 \$1960 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$38830 \$16 \$1860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38831 \$16 \$3461 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38832 \$16 \$1585 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38834 \$153 \$3534 \$3212 \$2192 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38835 \$16 \$3587 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38837 \$153 \$3568 \$3212 \$1860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38839 \$16 \$1960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38840 \$153 \$3440 \$3212 \$1960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38842 \$153 \$3534 \$2269 \$3167 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38843 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$38844 \$16 \$1960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38845 \$153 \$3568 \$2000 \$3167 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38846 \$153 \$3512 \$3250 \$1960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38847 \$16 \$4057 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38848 \$16 \$3373 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38849 \$153 \$3373 \$2192 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$38851 \$153 \$3512 \$2086 \$3342 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38852 \$153 \$3535 \$3250 \$2093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38853 \$16 \$2093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38854 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$38855 \$153 \$3535 \$2265 \$3342 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38856 \$153 \$3326 \$2267 \$3342 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38858 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$38859 \$16 \$1960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38860 \$16 \$2093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38861 \$153 \$3569 \$3147 \$1960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38862 \$153 \$3489 \$3147 \$2093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38863 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$38864 \$16 \$2085 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38865 \$153 \$3569 \$2086 \$3192 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38868 \$153 \$3489 \$2265 \$3192 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38869 \$16 \$3602 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38871 \$153 \$3265 \$2269 \$3192 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38872 \$16 \$1860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38873 \$153 \$3603 \$3251 \$1860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38874 \$153 \$3536 \$3251 \$2093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38876 \$153 \$3380 \$1936 \$3192 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38877 \$153 \$3441 \$3251 \$1960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38878 \$153 \$3536 \$2265 \$2931 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38880 \$153 \$3549 \$3252 \$2093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38881 \$16 \$2093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38882 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$38884 \$16 \$2085 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38885 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$38886 \$153 \$3549 \$2265 \$3169 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38888 \$153 \$3570 \$3252 \$1960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38889 \$16 \$1960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38891 \$16 \$1475 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38892 \$153 \$3469 \$2269 \$3169 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38894 \$16 \$2093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38896 \$153 \$3570 \$2086 \$3169 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38898 \$16 \$2093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38899 \$153 \$3442 \$3253 \$2093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38900 \$153 \$3443 \$3254 \$2093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38901 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$38904 \$16 \$3680 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38907 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$38908 \$16 \$1860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38909 \$16 \$1860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38910 \$153 \$3605 \$3254 \$1860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38911 \$153 \$3537 \$3253 \$1860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38912 \$153 \$3537 \$2000 \$3206 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38914 \$153 \$3538 \$3254 \$2192 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38916 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$38917 \$16 \$2192 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38918 \$153 \$3444 \$3253 \$2192 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38919 \$153 \$3539 \$3253 \$1960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38920 \$153 \$3539 \$2086 \$3206 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38921 \$16 \$1960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38923 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$38925 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$38926 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$38927 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$38928 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$38929 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$38930 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$38931 \$153 \$2286 \$3010 \$2006 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38932 \$153 \$2209 \$3010 \$1687 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38933 \$153 \$2287 \$3010 \$1658 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38934 \$16 \$2006 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38935 \$16 \$1687 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38936 \$16 \$1658 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38938 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$38939 \$153 \$2574 \$3010 \$2024 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38940 \$153 \$2687 \$1547 \$2785 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38941 \$153 \$2968 \$2009 \$2785 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38942 \$153 \$2669 \$3010 \$2180 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38945 \$153 \$3066 \$2064 \$2884 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38948 \$153 \$3207 \$1503 \$3137 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$38949 \$153 \$3067 \$2210 \$2884 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38951 \$16 \$981 \$2932 \$3037 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$38952 \$16 \$1496 \$2932 \$3137 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$38954 \$153 \$3092 \$2901 \$2024 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38956 \$153 \$3116 \$2901 \$2180 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38957 \$16 \$2024 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38958 \$16 \$2932 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38959 \$16 \$2180 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38960 \$153 \$3068 \$2064 \$3056 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38961 \$16 \$2932 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38962 \$16 \$1496 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38964 \$153 \$2849 \$2901 \$1942 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38967 \$153 \$3091 \$2009 \$2884 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38968 \$153 \$3116 \$2252 \$2886 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38969 \$153 \$3170 \$1686 \$3012 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$38970 \$153 \$3092 \$2210 \$2886 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38971 \$16 \$1404 \$16 \$153 \$3056 VNB sky130_fd_sc_hd__inv_1
X$38973 \$153 \$3069 \$2009 \$3056 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38976 \$153 \$3117 \$2887 \$1980 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38977 \$153 \$3013 \$2252 \$3014 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38978 \$153 \$2851 \$1792 \$3014 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38980 \$153 \$3070 \$3148 \$2180 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38983 \$153 \$3117 \$2009 \$3014 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38984 \$16 \$2180 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38985 \$16 \$1980 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38987 \$16 \$2932 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38988 \$16 \$1328 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38989 \$16 \$1328 \$2932 \$3057 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$38990 \$153 \$3171 \$3148 \$1687 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38991 \$153 \$3148 \$1576 \$3057 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$38993 \$16 \$1328 \$16 \$153 \$3149 VNB sky130_fd_sc_hd__inv_1
X$38994 \$153 \$3070 \$2252 \$3149 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$38995 \$16 \$1687 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38996 \$16 \$1328 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$38997 \$153 \$3016 \$3093 \$1687 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38998 \$153 \$3038 \$3093 \$2006 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$38999 \$153 \$3150 \$1547 \$3149 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39001 \$153 \$2810 \$2064 \$1594 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39003 \$153 \$2940 \$3093 \$1980 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39004 \$153 \$2763 \$1815 \$1594 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39005 \$16 \$1687 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39006 \$153 \$3093 \$1171 \$3039 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$39007 \$16 \$2442 \$16 \$153 \$2932 VNB sky130_fd_sc_hd__clkbuf_2
X$39008 \$16 \$1264 \$16 \$153 \$3015 VNB sky130_fd_sc_hd__inv_1
X$39010 \$16 \$2442 \$16 \$153 \$2647 VNB sky130_fd_sc_hd__clkbuf_2
X$39011 \$153 \$3118 \$3017 \$1658 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39012 \$153 \$2815 \$3017 \$2180 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39014 \$153 \$3119 \$3017 \$2006 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39015 \$16 \$2180 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39016 \$16 \$1658 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39017 \$16 \$2647 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39019 \$153 \$2837 \$3017 \$1980 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39020 \$16 \$1264 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39022 \$153 \$2591 \$3071 \$1795 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39023 \$16 \$1551 \$16 \$153 \$2743 VNB sky130_fd_sc_hd__inv_1
X$39024 \$153 \$3094 \$2933 \$1942 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39026 \$153 \$2672 \$3071 \$2024 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39027 \$153 \$2705 \$1547 \$2671 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39029 \$16 \$2180 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39030 \$16 \$1687 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39031 \$153 \$2975 \$1792 \$2889 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39032 \$16 \$1942 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39033 \$16 \$588 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39034 \$16 \$2006 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39035 \$153 \$2742 \$3071 \$2006 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39037 \$153 \$3040 \$3071 \$2180 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39039 \$16 \$2647 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39040 \$16 \$1354 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39041 \$16 \$2180 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39042 \$16 \$1658 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39043 \$153 \$3071 \$1332 \$3018 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$39044 \$153 \$153 \$2064 \$3151 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39046 \$153 \$3120 \$3071 \$1658 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39047 \$153 \$3095 \$3071 \$1980 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39048 \$153 \$153 \$2009 \$3151 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39049 \$16 \$1980 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39050 \$16 \$2878 \$16 \$153 \$1390 VNB sky130_fd_sc_hd__clkbuf_2
X$39051 \$16 \$1980 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39052 \$16 \$3490 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39054 \$153 \$3096 \$1980 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$39055 \$153 \$3019 \$2009 \$2889 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39057 \$153 \$3005 \$1503 \$3072 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$39058 \$153 \$2978 \$1895 \$2594 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39060 \$16 \$1923 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39061 \$153 \$3041 \$3020 \$1923 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39063 \$16 \$1547 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39064 \$16 \$2009 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39065 \$153 \$3073 \$3020 \$1965 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39067 \$153 \$3041 \$1895 \$3058 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39068 \$16 \$1965 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39070 \$153 \$3121 \$3020 \$2089 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39071 \$16 \$1923 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39074 \$153 \$3073 \$1806 \$3058 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39075 \$16 \$1923 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39076 \$153 \$3121 \$2026 \$3058 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39077 \$16 \$1503 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39078 \$153 \$2979 \$1954 \$2594 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39079 \$16 \$2089 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39080 \$153 \$3042 \$3020 \$2043 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39081 \$16 \$2042 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39082 \$16 \$981 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39083 \$16 \$1845 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39085 \$153 \$3074 \$3020 \$1805 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39086 \$153 \$3042 \$1954 \$3058 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39087 \$16 \$2043 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39089 \$153 \$3074 \$1703 \$3058 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39090 \$16 \$981 \$2539 \$3122 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$39091 \$153 \$3022 \$3144 \$1845 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39093 \$153 \$3144 \$1208 \$3122 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$39094 \$153 \$2859 \$3144 \$1805 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39095 \$153 \$3043 \$1924 \$2879 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39096 \$16 \$981 \$16 \$153 \$2879 VNB sky130_fd_sc_hd__inv_1
X$39097 \$153 \$3075 \$1806 \$2879 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39099 \$16 \$1805 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39100 \$16 \$1845 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39102 \$153 \$3153 \$1954 \$2879 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39103 \$153 \$3006 \$1686 \$3059 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$39104 \$153 \$3123 \$3006 \$2089 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39105 \$16 \$1404 \$2539 \$3059 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$39106 \$16 \$2539 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39108 \$16 \$1404 \$16 \$153 \$2925 VNB sky130_fd_sc_hd__inv_1
X$39109 \$153 \$3123 \$2026 \$2925 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39110 \$16 \$1404 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39111 \$16 \$1404 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39112 \$153 \$3044 \$3006 \$1923 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39113 \$153 \$3154 \$1806 \$2925 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39114 \$16 \$1576 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39115 \$16 \$2539 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39116 \$153 \$3044 \$1895 \$2925 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39117 \$16 \$2043 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39118 \$16 \$1923 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39120 \$153 \$3155 \$1703 \$2925 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39121 \$16 \$1328 \$2539 \$3045 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$39123 \$153 \$3097 \$2946 \$1923 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39125 \$153 \$3124 \$2946 \$2089 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39126 \$16 \$1923 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39127 \$16 \$2089 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39129 \$16 \$1328 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39130 \$16 \$1328 \$16 \$153 \$2895 VNB sky130_fd_sc_hd__inv_1
X$39131 \$16 \$3156 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39132 \$16 \$2199 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39133 \$16 \$3351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39134 \$16 \$1328 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39135 \$153 \$3125 \$2946 \$1965 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39136 \$153 \$2947 \$2946 \$1805 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39137 \$16 \$1965 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39138 \$16 \$1805 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39140 \$153 \$3023 \$1924 \$2895 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39141 \$16 \$1572 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39144 \$153 \$3157 \$1954 \$2895 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39145 \$16 \$2042 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39146 \$16 \$1171 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39147 \$16 \$2043 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39148 \$16 \$3240 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39149 \$153 \$3025 \$3024 \$2199 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39150 \$16 \$3352 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39152 \$153 \$3076 \$3024 \$2042 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39154 \$153 \$3076 \$1924 \$3060 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39155 \$16 \$1264 \$16 \$153 \$3060 VNB sky130_fd_sc_hd__inv_1
X$39156 \$16 \$2042 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39157 \$16 \$2199 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39158 \$153 \$2950 \$3024 \$1845 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39159 \$153 \$3026 \$3024 \$1805 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39160 \$16 \$1805 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39161 \$16 \$1845 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39162 \$16 \$1332 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39165 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$39166 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$39167 \$153 \$3126 \$3077 \$1923 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39168 \$153 \$3098 \$3077 \$1845 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39169 \$16 \$1923 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39170 \$16 \$1508 \$16 \$153 \$2908 VNB sky130_fd_sc_hd__inv_1
X$39171 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$39172 \$16 \$1845 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39173 \$153 \$3177 \$3077 \$2199 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39174 \$16 \$1508 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39177 \$153 \$3099 \$3077 \$1805 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39178 \$153 \$3158 \$2026 \$2908 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39179 \$16 \$1805 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39180 \$16 \$2908 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39182 \$16 \$2199 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39183 \$153 \$3046 \$2952 \$2042 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39185 \$16 \$1354 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39186 \$16 \$2908 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39188 \$153 \$3078 \$2952 \$2199 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39189 \$153 \$3046 \$1924 \$2926 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39190 \$153 \$3720 \$1805 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$39191 \$153 \$3078 \$2184 \$2926 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39193 \$153 \$3100 \$2952 \$2043 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39194 \$153 \$3100 \$1954 \$2926 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39195 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39196 \$153 \$3099 \$1703 \$2908 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39197 \$153 \$3047 \$1482 \$3354 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39198 \$16 \$3720 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39200 \$153 \$3096 \$1969 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$39201 \$153 \$2656 \$2863 \$1879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39202 \$153 \$3126 \$1895 \$2908 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39203 \$16 \$3079 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39205 \$16 \$3101 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39208 \$153 \$153 \$2438 \$3061 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39209 \$153 \$153 \$2092 \$3061 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39210 \$153 \$153 \$1558 \$3061 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39211 \$16 \$16 \$153 VNB sky130_fd_sc_hd__conb_1
X$39213 \$153 \$153 \$1868 \$3061 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39215 \$153 \$3027 \$2863 \$1878 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39216 \$16 \$1378 \$16 \$153 \$3061 VNB sky130_fd_sc_hd__clkbuf_2
X$39219 \$153 \$3127 \$3159 \$1989 \$3178 \$3145 \$2166 \$3139 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$39220 \$153 \$2997 \$1712 \$2639 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39222 \$16 \$1737 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39223 \$16 \$3272 \$3048 \$3081 \$1100 \$16 \$153 VNB sky130_fd_sc_hd__mux2_1
X$39225 \$153 \$3127 \$3128 \$1737 \$3047 \$3146 \$2774 \$3139 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$39227 \$153 \$3127 \$3138 \$1826 \$3102 \$3082 \$1650 \$3139 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$39228 \$153 \$3700 \$3788 \$3160 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39230 \$153 \$1368 \$21 \$1811 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39231 \$16 \$1969 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39232 \$16 \$1718 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39234 \$16 \$1879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39235 \$153 \$2998 \$1613 \$2752 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39236 \$153 \$3211 \$1933 \$2954 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$39237 \$153 \$3083 \$2696 \$2098 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39238 \$153 \$3129 \$2696 \$2105 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39241 \$153 \$3083 \$1993 \$2627 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39243 \$153 \$3163 \$1613 \$3162 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39244 \$153 \$3129 \$2438 \$2627 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39245 \$153 \$3282 \$1708 \$3104 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$39246 \$16 \$1518 \$2935 \$3104 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$39247 \$16 \$1756 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39248 \$153 \$3105 \$2796 \$1756 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39250 \$16 \$2659 \$16 \$153 \$2935 VNB sky130_fd_sc_hd__clkbuf_2
X$39251 \$153 \$3105 \$1712 \$2641 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39252 \$153 \$3140 \$1647 \$3106 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$39253 \$153 \$3062 \$1993 \$2641 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39254 \$16 \$1514 \$2935 \$3106 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$39256 \$153 \$3130 \$2866 \$2098 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39257 \$16 \$2098 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39259 \$16 \$2104 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39260 \$153 \$3029 \$2866 \$2104 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39261 \$153 \$3130 \$1993 \$2789 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39262 \$16 \$3048 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39263 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$39264 \$16 \$1514 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39265 \$16 \$1969 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39266 \$16 \$2016 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39268 \$153 \$3049 \$2866 \$2016 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39269 \$153 \$3180 \$2866 \$1969 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39270 \$153 \$3049 \$1715 \$2789 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39271 \$16 \$1758 \$2935 \$3181 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$39273 \$153 \$3007 \$2881 \$2105 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39274 \$16 \$2104 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39276 \$153 \$3107 \$2881 \$2104 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39277 \$16 \$1758 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39279 \$153 \$3107 \$2092 \$2790 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39280 \$16 \$2016 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39281 \$153 \$3050 \$2881 \$2016 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39282 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$39283 \$16 \$1599 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39285 \$153 \$3318 \$1558 \$3131 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39286 \$153 \$3050 \$1715 \$2790 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39287 \$16 \$1599 \$16 \$153 \$3131 VNB sky130_fd_sc_hd__inv_1
X$39288 \$153 \$3084 \$3085 \$2104 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39289 \$16 \$2104 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39290 \$16 \$1649 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39291 \$153 \$2868 \$1613 \$2791 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39293 \$153 \$3084 \$2092 \$3063 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39294 \$153 \$3182 \$3085 \$2098 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39295 \$153 \$3108 \$3085 \$2016 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39296 \$16 \$2016 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39298 \$153 \$3108 \$1715 \$3063 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39299 \$16 \$3087 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39300 \$16 \$2580 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39303 \$16 \$1228 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39304 \$16 \$2105 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39305 \$16 \$1121 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39306 \$153 \$3183 \$3085 \$2105 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39307 \$153 \$3085 \$1121 \$3051 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$39308 \$153 \$3132 \$3085 \$1756 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39310 \$16 \$1756 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39311 \$153 \$2983 \$1712 \$2791 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39312 \$153 \$3132 \$1712 \$3063 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39313 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39314 \$153 \$3109 \$1482 \$549 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39315 \$16 \$1228 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39317 \$16 \$3086 \$2960 \$3184 \$269 \$16 \$153 VNB sky130_fd_sc_hd__mux2_1
X$39319 \$16 \$549 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39320 \$153 \$3031 \$2958 \$2085 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39321 \$153 \$153 \$2056 \$3205 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39322 \$16 \$1044 \$16 \$153 \$2899 VNB sky130_fd_sc_hd__inv_1
X$39324 \$16 \$2085 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39325 \$153 \$153 \$2271 \$3205 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39326 \$153 \$153 \$2269 \$3205 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39327 \$16 \$2191 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39328 \$153 \$153 \$2000 \$3205 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39331 \$153 \$2871 \$2958 \$1973 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39332 \$16 \$1044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39333 \$16 \$1543 \$2984 \$3141 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$39334 \$153 \$3185 \$1760 \$3141 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$39335 \$153 \$3052 \$2958 \$1860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39337 \$16 \$1543 \$16 \$153 \$3186 VNB sky130_fd_sc_hd__inv_1
X$39338 \$16 \$2191 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39339 \$153 \$3052 \$2000 \$2899 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39340 \$16 \$1860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39342 \$153 \$3165 \$3142 \$3461 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39343 \$16 \$1585 \$2984 \$3110 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$39344 \$153 \$3089 \$2831 \$2085 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39345 \$153 \$3089 \$2271 \$2872 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39347 \$16 \$2085 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39348 \$153 \$2757 \$2000 \$2872 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39349 \$153 \$3212 \$1933 \$3110 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$39350 \$153 \$3053 \$2831 \$2192 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39351 \$153 \$3166 \$2056 \$3167 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39352 \$153 \$3053 \$2269 \$2872 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39354 \$16 \$2192 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39356 \$16 \$1960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39357 \$16 \$2191 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39359 \$153 \$3032 \$2832 \$2191 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39360 \$153 \$3189 \$2832 \$1960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39361 \$16 \$2803 \$16 \$153 \$2984 VNB sky130_fd_sc_hd__clkbuf_2
X$39362 \$16 \$1566 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39363 \$16 \$3064 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39365 \$16 \$3064 \$16 \$153 \$2803 VNB sky130_fd_sc_hd__clkbuf_2
X$39366 \$16 \$2085 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39367 \$16 \$2093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39368 \$153 \$3065 \$2832 \$2093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39369 \$153 \$3133 \$2832 \$2085 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39370 \$153 \$3065 \$2265 \$2780 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39371 \$16 \$1518 \$2984 \$3190 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$39372 \$16 \$2984 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39376 \$16 \$1518 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39377 \$16 \$1973 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39378 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$39379 \$153 \$3111 \$2874 \$1973 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39380 \$16 \$1973 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39381 \$153 \$3168 \$3147 \$1973 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39383 \$16 \$1514 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39385 \$16 \$2984 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39386 \$16 \$1860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39388 \$16 \$1514 \$2984 \$3193 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$39390 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$39391 \$153 \$3134 \$2874 \$1860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39393 \$16 \$2191 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39394 \$153 \$3054 \$2874 \$2191 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39395 \$153 \$3134 \$2000 \$2920 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39396 \$153 \$3054 \$2267 \$2920 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39399 \$16 \$1514 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39401 \$16 \$2085 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39402 \$16 \$1599 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39403 \$153 \$3112 \$2804 \$2085 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39404 \$16 \$1599 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39405 \$153 \$3194 \$2267 \$2931 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39406 \$16 \$1649 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39408 \$153 \$3112 \$2271 \$2759 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39409 \$16 \$1599 \$2984 \$3113 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$39412 \$153 \$2967 \$2804 \$1960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39413 \$16 \$1960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39415 \$16 \$1599 \$16 \$153 \$3169 VNB sky130_fd_sc_hd__inv_1
X$39416 \$16 \$1973 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39417 \$153 \$3195 \$2267 \$3169 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39418 \$153 \$3090 \$1121 \$2989 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$39419 \$153 \$3143 \$2271 \$2931 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39422 \$16 \$1758 \$2984 \$3196 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$39424 \$16 \$2093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39425 \$153 \$3114 \$3090 \$2093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39426 \$153 \$3135 \$3090 \$2085 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39427 \$16 \$1228 \$16 \$153 \$2923 VNB sky130_fd_sc_hd__inv_1
X$39428 \$153 \$3114 \$2265 \$2923 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39430 \$16 \$2191 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39432 \$153 \$3033 \$3090 \$2191 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39434 \$16 \$1860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39435 \$153 \$3034 \$3090 \$1860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39436 \$153 \$3115 \$3090 \$1973 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39437 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$39440 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$39442 \$16 \$1960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39443 \$16 \$2031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39444 \$153 \$3136 \$3090 \$1960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39445 \$153 \$3055 \$3090 \$2031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39446 \$153 \$3136 \$2086 \$2923 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39447 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$39450 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$39451 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$39452 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$39453 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$39454 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$39455 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$39457 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$39458 \$153 \$11362 \$11288 \$10427 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39460 \$153 \$11231 \$10276 \$11232 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39461 \$153 \$11286 \$10303 \$11232 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39462 \$16 \$10427 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39463 \$16 \$10368 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39464 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$39466 \$153 \$11287 \$10276 \$11263 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39468 \$153 \$11326 \$11288 \$10646 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39470 \$153 \$11189 \$11288 \$10367 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39471 \$153 \$11326 \$10318 \$11232 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39474 \$16 \$10367 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39475 \$16 \$11289 \$11347 \$11363 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$39477 \$16 \$11289 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39478 \$153 \$11264 \$11288 \$10476 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39479 \$153 \$11176 \$11288 \$10226 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39480 \$153 \$11264 \$10705 \$11232 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39481 \$16 \$11289 \$16 \$153 \$11232 VNB sky130_fd_sc_hd__inv_1
X$39482 \$16 \$10476 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39483 \$16 \$10226 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39485 \$153 \$11327 \$11348 \$10646 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39486 \$153 \$11233 \$11348 \$10368 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39487 \$153 \$11327 \$10318 \$11265 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39488 \$153 \$11233 \$10303 \$11265 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39489 \$16 \$10646 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39491 \$153 \$11328 \$11348 \$10367 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39493 \$153 \$11234 \$10705 \$10884 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39495 \$153 \$11235 \$10963 \$10200 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39496 \$153 \$11328 \$10330 \$11265 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39498 \$16 \$11274 \$16 \$153 \$10884 VNB sky130_fd_sc_hd__inv_1
X$39499 \$153 \$11235 \$10088 \$10884 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39502 \$153 \$10963 \$11190 \$11236 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$39503 \$16 \$10953 \$16 \$153 \$11347 VNB sky130_fd_sc_hd__clkbuf_2
X$39504 \$153 \$11192 \$11271 \$10295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39505 \$153 \$11193 \$11271 \$10368 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39507 \$153 \$11290 \$11271 \$10427 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39508 \$16 \$10427 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39509 \$16 \$10368 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39510 \$16 \$10295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39511 \$153 \$11290 \$10327 \$11191 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39513 \$153 \$11291 \$11271 \$10646 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39514 \$153 \$11468 \$10161 \$11191 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39517 \$16 \$10200 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39518 \$153 \$11291 \$10318 \$11191 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39519 \$153 \$11237 \$11271 \$10200 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39520 \$16 \$10646 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39521 \$16 \$10200 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39522 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$39523 \$153 \$11271 \$11364 \$11292 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$39524 \$16 \$10200 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39525 \$16 \$11297 \$10635 \$11292 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$39527 \$153 \$11237 \$10088 \$11191 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39528 \$16 \$11364 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39529 \$16 \$10427 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39530 \$153 \$11239 \$11000 \$10427 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39531 \$153 \$11365 \$11000 \$10226 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39532 \$16 \$10226 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39533 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$39536 \$153 \$11241 \$11000 \$10367 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39538 \$153 \$11178 \$11000 \$10200 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39539 \$153 \$11241 \$10330 \$10954 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39540 \$16 \$11240 \$16 \$153 \$10954 VNB sky130_fd_sc_hd__inv_1
X$39541 \$16 \$10476 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39542 \$153 \$11329 \$10971 \$10476 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39543 \$16 \$10367 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39546 \$16 \$11240 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39548 \$16 \$10427 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39549 \$153 \$11195 \$10971 \$10427 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39550 \$153 \$11329 \$10705 \$11057 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39551 \$153 \$11158 \$10161 \$11057 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39552 \$153 \$11293 \$10971 \$10200 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39554 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$39555 \$153 \$10971 \$11431 \$11338 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$39556 \$153 \$11293 \$10088 \$11057 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39557 \$16 \$10974 \$11238 \$11242 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$39558 \$16 \$11267 \$11238 \$11338 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$39559 \$16 \$11266 \$16 \$153 \$10555 VNB sky130_fd_sc_hd__clkbuf_2
X$39560 \$16 \$11431 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39561 \$16 \$11349 \$16 \$153 \$11297 VNB sky130_fd_sc_hd__clkbuf_2
X$39563 \$16 \$11267 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39564 \$153 \$11349 \$11197 \$11159 \$11243 \$11180 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$39565 \$153 \$11266 \$11197 \$11243 \$11180 \$11159 \$16 \$16 VNB
+ sky130_fd_sc_hd__nor4b_2
X$39566 \$153 \$11243 \$11197 \$11350 \$11180 \$11159 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$39567 \$153 \$11118 \$11180 \$11159 \$11243 \$11197 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$39568 \$16 \$11295 \$16 \$153 \$10413 VNB sky130_fd_sc_hd__clkbuf_2
X$39569 \$153 \$11197 \$11180 \$11294 \$11243 \$11159 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$39570 \$16 \$11244 \$16 \$153 \$11243 VNB sky130_fd_sc_hd__clkbuf_2
X$39572 \$153 \$11243 \$11180 \$11352 \$11197 \$11159 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$39573 \$16 \$11159 \$11180 \$11243 \$11197 \$16 \$153 \$11295 VNB
+ sky130_fd_sc_hd__and4_2
X$39575 \$16 \$11272 \$11273 \$11296 \$153 \$16 \$11351 VNB
+ sky130_fd_sc_hd__and3_4
X$39576 \$16 \$11119 \$16 \$153 \$11197 VNB sky130_fd_sc_hd__clkbuf_2
X$39578 \$16 \$11273 \$11296 \$11272 \$153 \$11198 \$16 VNB
+ sky130_fd_sc_hd__and3b_4
X$39579 \$153 \$11273 \$11272 \$11366 \$11296 \$16 \$16 VNB
+ sky130_fd_sc_hd__nor3b_4
X$39581 \$16 \$7801 \$16 \$153 \$11273 VNB sky130_fd_sc_hd__clkbuf_2
X$39582 \$16 \$7656 \$16 \$153 \$11272 VNB sky130_fd_sc_hd__clkbuf_2
X$39583 \$16 \$10500 \$16 \$153 \$11296 VNB sky130_fd_sc_hd__clkbuf_2
X$39584 \$16 \$7801 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39585 \$16 \$10500 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39587 \$153 \$11298 \$11120 \$10514 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39588 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$39589 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$39590 \$16 \$10526 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39592 \$16 \$10514 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39593 \$16 \$11289 \$16 \$153 \$11200 VNB sky130_fd_sc_hd__inv_1
X$39594 \$153 \$11137 \$10344 \$11200 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39595 \$16 \$10605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39596 \$16 \$11289 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39597 \$153 \$11367 \$11120 \$10338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39598 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$39599 \$153 \$11368 \$11120 \$10470 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39600 \$16 \$10338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39601 \$16 \$11274 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39603 \$153 \$11182 \$11120 \$10382 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39604 \$153 \$11121 \$11190 \$11339 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$39605 \$16 \$11274 \$11275 \$11339 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$39606 \$153 \$11122 \$11121 \$10298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39607 \$16 \$10382 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39610 \$16 \$10470 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39611 \$16 \$11190 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39612 \$16 \$11567 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39613 \$16 \$11369 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39614 \$153 \$11370 \$10344 \$11112 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39616 \$153 \$11245 \$10309 \$11112 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39617 \$16 \$10298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39618 \$153 \$11138 \$10098 \$11112 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39619 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$39620 \$153 \$11340 \$10247 \$11112 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39622 \$153 \$11341 \$11121 \$10526 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39623 \$153 \$11341 \$10516 \$11112 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39624 \$16 \$11274 \$16 \$153 \$11112 VNB sky130_fd_sc_hd__inv_1
X$39625 \$153 \$11299 \$11060 \$10338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39627 \$153 \$11299 \$10309 \$10956 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39629 \$16 \$11274 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39630 \$153 \$11183 \$11060 \$10605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39631 \$153 \$11201 \$11060 \$10606 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39632 \$16 \$10605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39633 \$16 \$10606 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39634 \$16 \$11364 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39635 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$39636 \$153 \$11124 \$11364 \$11342 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$39638 \$16 \$11297 \$10655 \$11342 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$39639 \$16 \$11297 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39641 \$153 \$11202 \$11124 \$10514 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39642 \$153 \$11184 \$11124 \$10526 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39643 \$16 \$10514 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39644 \$16 \$10526 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39646 \$16 \$11297 \$16 \$153 \$10958 VNB sky130_fd_sc_hd__inv_1
X$39649 \$16 \$11297 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39650 \$153 \$11203 \$11124 \$10605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39651 \$153 \$11246 \$11124 \$10382 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39652 \$153 \$11246 \$10098 \$10958 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39653 \$16 \$10382 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39654 \$16 \$6328 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39655 \$16 \$6328 \$16 \$153 \$7894 VNB sky130_fd_sc_hd__clkbuf_2
X$39656 \$153 \$11049 \$11194 \$11301 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$39658 \$153 \$11300 \$11049 \$10338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39659 \$16 \$11077 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39660 \$153 \$11300 \$10309 \$11061 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39661 \$16 \$11077 \$10655 \$11301 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$39663 \$153 \$11302 \$11049 \$10382 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39664 \$16 \$11077 \$16 \$153 \$11061 VNB sky130_fd_sc_hd__inv_1
X$39665 \$16 \$10382 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39667 \$153 \$11303 \$11049 \$10470 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39668 \$16 \$10382 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39669 \$153 \$11247 \$11276 \$10470 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39670 \$16 \$10470 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39671 \$153 \$11371 \$11276 \$10298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39673 \$153 \$11303 \$10247 \$11061 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39674 \$16 \$10338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39675 \$153 \$11277 \$11276 \$10605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39676 \$16 \$10974 \$11164 \$11206 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$39677 \$153 \$11304 \$11276 \$10382 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39678 \$16 \$10298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39679 \$16 \$10298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39681 \$153 \$11304 \$10098 \$11205 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39682 \$153 \$11277 \$10686 \$11205 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39683 \$16 \$11267 \$11164 \$11372 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$39685 \$153 \$11305 \$11208 \$10298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39686 \$16 \$10514 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39687 \$153 \$11330 \$11208 \$10514 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39689 \$16 \$11267 \$16 \$153 \$11268 VNB sky130_fd_sc_hd__inv_1
X$39690 \$153 \$11330 \$10538 \$11268 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39691 \$153 \$11305 \$10401 \$11268 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39692 \$16 \$10605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39693 \$153 \$11373 \$10098 \$11906 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39694 \$16 \$11267 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39696 \$16 \$10526 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39697 \$153 \$11249 \$11208 \$10526 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39698 \$16 \$11267 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39699 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$39701 \$16 \$10470 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39703 \$153 \$11353 \$10247 \$11268 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39704 \$153 \$11249 \$10516 \$11268 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39706 \$16 \$10735 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39707 \$153 \$11142 \$10686 \$10894 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39708 \$153 \$11331 \$11050 \$10735 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39709 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$39711 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$39712 \$153 \$11331 \$10919 \$11209 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39714 \$153 \$11210 \$11050 \$10578 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39715 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$39716 \$153 \$11306 \$11050 \$10551 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39717 \$16 \$10578 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39719 \$16 \$11374 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39721 \$16 \$11374 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39722 \$16 \$11113 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39723 \$153 \$11306 \$10471 \$11209 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39725 \$153 \$11050 \$11148 \$11250 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$39726 \$16 \$11113 \$16 \$153 \$11209 VNB sky130_fd_sc_hd__inv_1
X$39728 \$16 \$10735 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39729 \$153 \$11332 \$11185 \$10735 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39730 \$16 \$10551 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39731 \$16 \$10735 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39732 \$16 \$10386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39734 \$16 \$11148 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39735 \$16 \$11113 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39736 \$16 \$11207 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39737 \$16 \$10809 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39738 \$153 \$11375 \$11185 \$10473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39739 \$153 \$11251 \$11185 \$10809 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39740 \$16 \$10473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39741 \$153 \$11251 \$10714 \$11065 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39743 \$16 \$10611 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39745 \$153 \$11332 \$10919 \$11065 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39747 \$153 \$11211 \$10979 \$10551 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39748 \$153 \$11377 \$11410 \$10611 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39749 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$39750 \$153 \$11376 \$10472 \$11354 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39751 \$16 \$10473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39754 \$153 \$11307 \$10979 \$10473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39756 \$153 \$10979 \$12347 \$11308 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$39757 \$16 \$11013 \$11127 \$11308 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$39758 \$16 \$11212 \$16 \$153 \$11378 VNB sky130_fd_sc_hd__clkbuf_2
X$39759 \$16 \$11013 \$16 \$153 \$10810 VNB sky130_fd_sc_hd__inv_1
X$39761 \$153 \$11252 \$10881 \$10300 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39762 \$16 \$10386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39764 \$153 \$11213 \$10881 \$10386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39765 \$153 \$11252 \$10417 \$10946 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39766 \$153 \$11307 \$10501 \$10810 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39768 \$16 \$11214 \$11378 \$11269 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$39769 \$153 \$11333 \$11355 \$10611 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39771 \$153 \$10881 \$11216 \$11269 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$39772 \$153 \$11379 \$10472 \$11215 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39773 \$16 \$10611 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39775 \$16 \$10473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39776 \$153 \$11309 \$11355 \$10473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39777 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$39779 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$39780 \$153 \$11356 \$10919 \$11215 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39782 \$16 \$11212 \$16 \$153 \$11412 VNB sky130_fd_sc_hd__clkbuf_2
X$39783 \$153 \$11217 \$11278 \$10809 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39785 \$16 \$10735 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39786 \$153 \$11380 \$11278 \$10735 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39788 \$153 \$10405 \$10472 \$10757 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39789 \$16 \$10661 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39790 \$16 \$10611 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39791 \$16 \$10473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39792 \$153 \$11130 \$11278 \$10473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39793 \$153 \$10983 \$11278 \$10611 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39794 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$39795 \$16 \$10552 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39796 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$39799 \$16 \$10551 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39800 \$16 \$10735 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39801 \$153 \$11218 \$11279 \$10551 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39802 \$153 \$11187 \$11279 \$10735 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39804 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$39805 \$16 \$10473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39806 \$153 \$11220 \$11279 \$10473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39807 \$16 \$10578 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39809 \$153 \$11310 \$11279 \$10578 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39810 \$153 \$11310 \$10370 \$11219 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39812 \$16 \$10611 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39813 \$153 \$11343 \$10472 \$11270 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39814 \$16 \$10473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39815 \$153 \$11131 \$11066 \$10611 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39817 \$153 \$11343 \$11311 \$10386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39818 \$153 \$11334 \$11311 \$10473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39819 \$16 \$10386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39820 \$16 \$11172 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39821 \$16 \$10300 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39822 \$16 \$10551 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39824 \$153 \$11312 \$11311 \$10300 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39825 \$16 \$10809 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39827 \$153 \$11344 \$11311 \$10809 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39828 \$153 \$11344 \$10714 \$11270 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39829 \$16 \$11412 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39830 \$153 \$11066 \$11280 \$11313 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$39831 \$16 \$11172 \$11412 \$11313 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$39832 \$16 \$7801 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39834 \$16 \$7801 \$16 \$153 \$11357 VNB sky130_fd_sc_hd__clkbuf_2
X$39835 \$153 \$11312 \$10417 \$11270 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39836 \$16 \$11359 \$11358 \$11357 \$153 \$11221 \$16 VNB
+ sky130_fd_sc_hd__and3b_4
X$39837 \$16 \$10986 \$16 \$153 \$11254 VNB sky130_fd_sc_hd__clkbuf_2
X$39838 \$16 \$7559 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39839 \$153 \$11133 \$11222 \$11223 \$11255 \$11254 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$39841 \$153 \$11381 \$11255 \$11223 \$11222 \$11254 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$39844 \$153 \$11382 \$11222 \$11255 \$11254 \$11223 \$16 \$16 VNB
+ sky130_fd_sc_hd__nor4b_2
X$39846 \$16 \$11016 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39847 \$153 \$11255 \$11222 \$11314 \$11254 \$11223 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$39848 \$16 \$11223 \$11254 \$11255 \$11222 \$16 \$153 \$11383 VNB
+ sky130_fd_sc_hd__and4_2
X$39849 \$153 \$11222 \$11254 \$10989 \$11255 \$11223 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$39850 \$153 \$11360 \$10642 \$11016 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39851 \$153 \$11345 \$11281 \$10564 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39853 \$16 \$11314 \$16 \$153 \$10831 VNB sky130_fd_sc_hd__clkbuf_2
X$39854 \$153 \$11345 \$10642 \$11226 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39856 \$16 \$10564 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39857 \$153 \$11225 \$11281 \$10326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39858 \$153 \$11315 \$11281 \$10467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39861 \$16 \$10467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39862 \$153 \$11315 \$10587 \$11226 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39863 \$16 \$10326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39865 \$153 \$11282 \$11281 \$10346 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39866 \$16 \$11113 \$16 \$153 \$10961 VNB sky130_fd_sc_hd__inv_1
X$39867 \$153 \$11282 \$10285 \$11226 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39868 \$153 \$11256 \$11281 \$10393 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39869 \$16 \$10346 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39870 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$39872 \$153 \$11335 \$11281 \$10446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39873 \$153 \$11256 \$10694 \$11226 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39874 \$153 \$11335 \$10376 \$11226 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39875 \$153 \$11257 \$10376 \$10961 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39876 \$153 \$11336 \$11316 \$10346 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39878 \$16 \$11013 \$10838 \$11258 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$39879 \$16 \$10564 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39880 \$153 \$11336 \$10285 \$11384 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39881 \$153 \$11361 \$10694 \$11384 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39882 \$153 \$11317 \$11316 \$10564 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39883 \$16 \$10346 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39884 \$16 \$10446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39885 \$16 \$10326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39887 \$16 \$10392 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39888 \$153 \$11317 \$10642 \$11384 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39890 \$16 \$10326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39891 \$16 \$11214 \$11504 \$11259 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$39892 \$16 \$11214 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39893 \$153 \$11228 \$11283 \$10326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39894 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$39895 \$153 \$11284 \$11283 \$10346 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39897 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$39898 \$153 \$11284 \$10285 \$11495 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39899 \$16 \$10346 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39901 \$16 \$10392 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39902 \$16 \$10393 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39903 \$153 \$11260 \$11283 \$10393 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39904 \$153 \$11337 \$11283 \$10392 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39906 \$153 \$11260 \$10694 \$11495 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39907 \$153 \$11337 \$10815 \$11495 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39909 \$16 \$10346 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39910 \$16 \$10467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39911 \$153 \$10486 \$11346 \$10346 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39912 \$153 \$11102 \$11346 \$10326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39913 \$16 \$10326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39915 \$16 \$10990 \$16 \$153 \$11229 VNB sky130_fd_sc_hd__clkbuf_2
X$39916 \$16 \$10392 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39917 \$16 \$10393 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39919 \$153 \$11068 \$11346 \$10392 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39920 \$153 \$11318 \$11346 \$10393 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39922 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$39923 \$16 \$11385 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39924 \$16 \$11280 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39926 \$16 \$10346 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39927 \$16 \$10326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39929 \$153 \$11319 \$11285 \$10346 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39930 \$153 \$11386 \$11285 \$10326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39931 \$16 \$10617 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39933 \$153 \$10364 \$10466 \$10650 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39934 \$153 \$11391 \$11285 \$10617 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39937 \$153 \$11320 \$11285 \$10392 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39938 \$153 \$11107 \$10560 \$11516 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39939 \$153 \$11053 \$11280 \$11262 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$39941 \$153 \$11321 \$11053 \$10564 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39943 \$153 \$10798 \$10285 \$11022 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39944 \$16 \$11172 \$16 \$153 \$11322 VNB sky130_fd_sc_hd__inv_1
X$39945 \$153 \$11323 \$11053 \$10617 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39946 \$153 \$10568 \$10560 \$10801 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39947 \$153 \$11387 \$11230 \$10393 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39948 \$16 \$10393 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39949 \$16 \$10326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39951 \$153 \$10936 \$10694 \$11022 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39952 \$153 \$11589 \$11230 \$10346 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39953 \$153 \$11324 \$11230 \$10326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39954 \$16 \$10346 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39955 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$39956 \$153 \$10802 \$10466 \$10741 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39959 \$16 \$10467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39960 \$153 \$11388 \$11230 \$10467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39961 \$153 \$11325 \$11230 \$10446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39962 \$153 \$10804 \$10560 \$10741 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39963 \$16 \$10510 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39964 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$39966 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$39967 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$39969 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$39970 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$39971 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$39972 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$39975 \$153 \$11518 \$11499 \$10427 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39976 \$153 \$11287 \$11499 \$10295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39977 \$153 \$11518 \$10327 \$11263 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39978 \$16 \$10295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39979 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$39980 \$16 \$10427 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39982 \$153 \$11519 \$10303 \$11263 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39983 \$153 \$11521 \$11499 \$10646 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39984 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$39986 \$153 \$11520 \$10088 \$11263 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39987 \$153 \$11521 \$10318 \$11263 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39988 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$39991 \$16 \$10646 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39992 \$153 \$11499 \$11720 \$11630 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$39993 \$16 \$11636 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39994 \$16 \$11636 \$16 \$153 \$11263 VNB sky130_fd_sc_hd__inv_1
X$39995 \$153 \$11591 \$11499 \$10226 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$39996 \$16 \$11636 \$11347 \$11630 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$39997 \$153 \$11591 \$10161 \$11263 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$39998 \$16 \$10226 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$39999 \$16 \$11636 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40000 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$40002 \$16 \$11720 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40003 \$153 \$11522 \$11348 \$10226 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40004 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$40005 \$153 \$11684 \$11751 \$10646 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40006 \$153 \$11522 \$10161 \$11265 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40007 \$16 \$10476 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40008 \$16 \$10646 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40009 \$16 \$10295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40011 \$153 \$11685 \$11631 \$10476 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40013 \$16 \$10226 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40014 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$40015 \$16 \$11369 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40016 \$153 \$11348 \$11567 \$11523 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$40017 \$153 \$11649 \$10276 \$11650 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40018 \$16 \$11567 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40019 \$16 \$11369 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40020 \$16 \$10476 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40021 \$153 \$11592 \$11631 \$10646 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40022 \$16 \$10427 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40024 \$153 \$11686 \$11631 \$10427 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40025 \$153 \$11592 \$10318 \$11650 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40026 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$40027 \$16 \$10646 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40028 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$40029 \$153 \$11614 \$11632 \$10646 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40031 \$16 \$10367 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40032 \$16 \$10427 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40033 \$153 \$11568 \$10276 \$11560 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40034 \$153 \$11614 \$10318 \$11560 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40035 \$153 \$11423 \$11484 \$10427 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40036 \$16 \$10646 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40037 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$40041 \$153 \$11177 \$11484 \$10295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40042 \$153 \$11469 \$11633 \$10295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40043 \$153 \$11524 \$10303 \$11393 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40044 \$153 \$11401 \$11484 \$10226 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40045 \$16 \$10295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40047 \$16 \$10295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40048 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$40049 \$16 \$10226 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40050 \$153 \$11651 \$10327 \$11652 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40051 \$153 \$11525 \$10318 \$11393 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40052 \$153 \$11634 \$10318 \$11652 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40053 \$153 \$11593 \$11484 \$10367 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40054 \$16 \$10476 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40055 \$16 \$11485 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40057 \$153 \$11615 \$10088 \$11652 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40058 \$153 \$11593 \$10330 \$11393 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40059 \$16 \$10367 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40060 \$153 \$11569 \$11735 \$10295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40061 \$16 \$11485 \$16 \$153 \$11393 VNB sky130_fd_sc_hd__inv_1
X$40063 \$16 \$10367 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40064 \$153 \$11569 \$10276 \$11719 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40065 \$153 \$11402 \$11425 \$10476 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40067 \$153 \$11505 \$11425 \$10367 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40068 \$153 \$11653 \$10318 \$11719 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40069 \$16 \$11485 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40070 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$40072 \$153 \$11595 \$11425 \$10295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40074 \$16 \$11594 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40076 \$16 \$10295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40077 \$16 \$11594 \$11238 \$11635 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$40078 \$153 \$11425 \$11689 \$11635 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$40080 \$153 \$11526 \$11425 \$10200 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40081 \$16 \$11689 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40083 \$16 \$11594 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40084 \$16 \$11594 \$16 \$153 \$11395 VNB sky130_fd_sc_hd__inv_1
X$40086 \$153 \$11526 \$10088 \$11395 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40087 \$16 \$10646 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40088 \$16 \$10200 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40089 \$153 \$11654 \$10276 \$11655 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40090 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$40092 \$16 \$11527 \$16 \$153 \$11240 VNB sky130_fd_sc_hd__clkbuf_2
X$40093 \$16 \$11814 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40095 \$153 \$11570 \$11428 \$11427 \$11429 \$11430 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$40096 \$16 \$11570 \$16 \$153 \$11485 VNB sky130_fd_sc_hd__clkbuf_2
X$40098 \$16 \$11506 \$16 \$153 \$11267 VNB sky130_fd_sc_hd__clkbuf_2
X$40099 \$153 \$11429 \$11430 \$11596 \$11428 \$11427 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$40101 \$153 \$11428 \$11430 \$11690 \$11429 \$11427 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$40103 \$16 \$11596 \$16 \$153 \$10974 VNB sky130_fd_sc_hd__clkbuf_2
X$40104 \$16 \$11111 \$16 \$153 \$11561 VNB sky130_fd_sc_hd__clkbuf_2
X$40105 \$16 \$11572 \$16 \$153 \$11369 VNB sky130_fd_sc_hd__clkbuf_2
X$40107 \$153 \$11571 \$11507 \$11508 \$11561 \$11529 \$16 \$16 VNB
+ sky130_fd_sc_hd__nor4b_2
X$40108 \$16 \$11528 \$16 \$153 \$11289 VNB sky130_fd_sc_hd__clkbuf_2
X$40109 \$16 \$11571 \$16 \$153 \$11274 VNB sky130_fd_sc_hd__clkbuf_2
X$40111 \$153 \$11500 \$11720 \$11691 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$40113 \$153 \$11572 \$11508 \$11529 \$11507 \$11561 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$40114 \$16 \$11366 \$16 \$153 \$11529 VNB sky130_fd_sc_hd__clkbuf_2
X$40115 \$153 \$11616 \$11500 \$10514 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40116 \$153 \$11434 \$11500 \$10605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40119 \$153 \$11530 \$10516 \$11396 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40120 \$153 \$11616 \$10538 \$11396 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40121 \$16 \$10605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40122 \$153 \$11656 \$10344 \$11396 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40124 \$153 \$11487 \$10309 \$11396 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40125 \$16 \$11636 \$16 \$153 \$11396 VNB sky130_fd_sc_hd__inv_1
X$40126 \$16 \$11636 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40127 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$40128 \$153 \$11617 \$11500 \$10382 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40130 \$153 \$11531 \$11500 \$10298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40131 \$153 \$11617 \$10098 \$11396 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40132 \$153 \$11531 \$10401 \$11396 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40133 \$16 \$10298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40134 \$16 \$10382 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40137 \$153 \$11435 \$11567 \$11532 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$40138 \$16 \$10470 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40140 \$153 \$11618 \$11657 \$10470 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40141 \$153 \$11597 \$11435 \$10470 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40142 \$153 \$11619 \$11657 \$10382 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40144 \$16 \$11369 \$16 \$153 \$11397 VNB sky130_fd_sc_hd__inv_1
X$40145 \$153 \$11533 \$10401 \$11397 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40146 \$153 \$11597 \$10247 \$11397 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40147 \$16 \$10470 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40148 \$16 \$10382 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40149 \$16 \$10470 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40150 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$40152 \$153 \$11509 \$11435 \$10338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40156 \$153 \$11573 \$11658 \$10470 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40157 \$153 \$11436 \$10686 \$11397 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40158 \$16 \$10338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40160 \$153 \$11573 \$10247 \$11562 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40161 \$153 \$11659 \$10401 \$11562 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40162 \$16 \$11485 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40163 \$16 \$10470 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40165 \$153 \$11534 \$10516 \$11397 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40167 \$16 \$11637 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40168 \$153 \$11661 \$10309 \$11660 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40169 \$153 \$11474 \$10538 \$11397 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40170 \$153 \$11439 \$11637 \$11694 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$40171 \$153 \$11406 \$11439 \$10470 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40172 \$16 \$11164 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40174 \$153 \$11662 \$10247 \$11660 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40175 \$153 \$11598 \$11439 \$10605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40176 \$153 \$11638 \$10098 \$11660 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40177 \$153 \$11598 \$10686 \$11398 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40178 \$16 \$11485 \$16 \$153 \$11398 VNB sky130_fd_sc_hd__inv_1
X$40179 \$16 \$10470 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40182 \$16 \$10605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40183 \$153 \$11599 \$11439 \$10298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40184 \$153 \$11663 \$10309 \$11488 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40185 \$153 \$11695 \$11639 \$10382 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40186 \$153 \$11600 \$11439 \$10606 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40187 \$16 \$10298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40189 \$153 \$11599 \$10401 \$11398 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40190 \$16 \$10298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40191 \$16 \$10382 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40192 \$153 \$11276 \$11856 \$11535 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$40193 \$16 \$10338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40194 \$16 \$10606 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40195 \$16 \$11795 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40196 \$16 \$11164 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40197 \$153 \$11407 \$11276 \$10606 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40198 \$16 \$11856 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40199 \$16 \$11689 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40200 \$16 \$11795 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40202 \$153 \$11574 \$10247 \$11563 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40203 \$153 \$11664 \$10401 \$11563 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40204 \$16 \$11240 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40206 \$16 \$11164 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40207 \$16 \$10606 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40208 \$153 \$11510 \$11276 \$10514 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40209 \$16 \$10606 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40210 \$153 \$11640 \$10098 \$11563 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40213 \$16 \$10514 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40214 \$153 \$11536 \$10309 \$11205 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40215 \$153 \$11696 \$11575 \$10606 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40217 \$153 \$11601 \$11575 \$10382 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40218 \$153 \$11620 \$11575 \$10514 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40220 \$153 \$11576 \$10401 \$11564 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40221 \$153 \$11620 \$10538 \$11564 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40222 \$16 \$11488 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40224 \$16 \$10338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40225 \$153 \$11537 \$11575 \$10338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40226 \$153 \$11696 \$10344 \$11564 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40227 \$16 \$10470 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40228 \$16 \$10526 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40230 \$153 \$11697 \$11575 \$10526 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40231 \$153 \$11602 \$11575 \$10470 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40232 \$16 \$11594 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40233 \$153 \$11537 \$10309 \$11564 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40234 \$16 \$10735 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40236 \$16 \$10809 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40237 \$153 \$11698 \$11501 \$10809 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40240 \$153 \$11603 \$11501 \$10300 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40242 \$153 \$11408 \$11501 \$10551 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40244 \$153 \$10829 \$11501 \$10611 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40246 \$16 \$10551 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40248 \$153 \$11501 \$11451 \$11538 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$40249 \$16 \$11374 \$16 \$153 \$11207 VNB sky130_fd_sc_hd__inv_1
X$40250 \$16 \$11399 \$11127 \$11577 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$40251 \$153 \$11185 \$11578 \$11577 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$40252 \$153 \$11621 \$11641 \$10611 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40255 \$153 \$11409 \$11185 \$10551 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40256 \$153 \$11797 \$10714 \$11665 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40257 \$153 \$11621 \$10833 \$11665 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40258 \$153 \$11512 \$11185 \$10300 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40259 \$16 \$10611 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40261 \$16 \$10386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40263 \$153 \$11700 \$11666 \$10386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40264 \$16 \$11578 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40266 \$16 \$10473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40267 \$153 \$11539 \$11410 \$10473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40268 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$40269 \$153 \$11377 \$10833 \$11354 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40270 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$40272 \$153 \$11539 \$10501 \$11354 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40273 \$153 \$11667 \$10919 \$11513 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40274 \$153 \$11579 \$10370 \$11513 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40275 \$16 \$10551 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40276 \$16 \$10611 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40278 \$153 \$11642 \$10714 \$11354 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40279 \$153 \$11540 \$10471 \$11354 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40282 \$153 \$11668 \$10833 \$11669 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40284 \$16 \$11502 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40285 \$16 \$11502 \$11378 \$11565 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$40286 \$153 \$11410 \$11604 \$11565 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$40287 \$153 \$11541 \$10370 \$11354 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40288 \$153 \$11643 \$10501 \$11669 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40289 \$16 \$11604 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40291 \$16 \$10300 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40293 \$153 \$11355 \$12612 \$11670 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$40294 \$153 \$11644 \$11355 \$10300 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40295 \$153 \$11644 \$10417 \$11215 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40296 \$16 \$10578 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40297 \$153 \$11605 \$11355 \$10578 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40298 \$16 \$12612 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40300 \$16 \$11622 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40302 \$16 \$11622 \$16 \$153 \$11215 VNB sky130_fd_sc_hd__inv_1
X$40303 \$153 \$11605 \$10370 \$11215 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40304 \$153 \$11514 \$11355 \$10809 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40306 \$16 \$10386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40307 \$153 \$11623 \$11278 \$10386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40308 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$40310 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$40311 \$153 \$11446 \$10417 \$10948 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40312 \$153 \$11542 \$10471 \$10948 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40313 \$153 \$11623 \$10472 \$10948 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40314 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$40315 \$16 \$11585 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40316 \$153 \$11278 \$11585 \$11543 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$40318 \$16 \$11627 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40319 \$16 \$10611 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40320 \$16 \$10300 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40322 \$153 \$11624 \$11645 \$10611 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40324 \$153 \$11448 \$11279 \$10300 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40325 \$153 \$11671 \$10501 \$11727 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40327 \$16 \$11413 \$16 \$153 \$11219 VNB sky130_fd_sc_hd__inv_1
X$40329 \$16 \$11413 \$11412 \$11672 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$40331 \$153 \$11544 \$10714 \$11219 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40332 \$153 \$11279 \$12404 \$11672 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$40333 \$153 \$11545 \$10833 \$11219 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40334 \$16 \$10578 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40335 \$153 \$11606 \$11580 \$10578 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40336 \$153 \$11674 \$10833 \$11673 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40338 \$16 \$12404 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40340 \$16 \$10473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40341 \$16 \$11413 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40342 \$153 \$11414 \$11580 \$10473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40343 \$153 \$11606 \$10370 \$11673 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40344 \$153 \$11701 \$10472 \$11673 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40345 \$16 \$10735 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40347 \$16 \$11546 \$16 \$153 \$11270 VNB sky130_fd_sc_hd__inv_1
X$40349 \$16 \$10809 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40351 \$153 \$11625 \$11580 \$10300 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40352 \$153 \$11547 \$10833 \$11270 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40353 \$16 \$10551 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40354 \$153 \$11548 \$11580 \$10551 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40356 \$153 \$11625 \$10417 \$11673 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40357 \$16 \$11280 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40358 \$153 \$11548 \$10471 \$11673 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40360 \$16 \$11459 \$16 \$153 \$11673 VNB sky130_fd_sc_hd__inv_1
X$40362 \$16 \$11675 \$16 \$153 \$11459 VNB sky130_fd_sc_hd__clkbuf_2
X$40363 \$16 \$11412 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40364 \$16 \$11676 \$16 \$153 \$11413 VNB sky130_fd_sc_hd__clkbuf_2
X$40366 \$16 \$11359 \$11357 \$11358 \$153 \$16 \$11581 VNB
+ sky130_fd_sc_hd__and3_4
X$40367 \$16 \$10986 \$16 \$153 \$11646 VNB sky130_fd_sc_hd__clkbuf_2
X$40368 \$16 \$11253 \$16 \$153 \$11626 VNB sky130_fd_sc_hd__clkbuf_2
X$40369 \$16 \$11549 \$16 \$153 \$11803 VNB sky130_fd_sc_hd__clkbuf_2
X$40370 \$153 \$11676 \$11582 \$11607 \$11626 \$11646 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$40371 \$16 \$11581 \$16 \$153 \$11607 VNB sky130_fd_sc_hd__clkbuf_2
X$40374 \$16 \$11578 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40375 \$153 \$11675 \$11626 \$11607 \$11582 \$11646 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$40376 \$16 \$11374 \$10838 \$11416 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$40377 \$153 \$11626 \$11646 \$11608 \$11582 \$11607 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$40378 \$16 \$11224 \$16 \$153 \$10739 VNB sky130_fd_sc_hd__clkbuf_2
X$40379 \$16 \$11374 \$16 \$153 \$11515 VNB sky130_fd_sc_hd__inv_1
X$40380 \$153 \$11609 \$11452 \$10392 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40381 \$153 \$11647 \$10466 \$11515 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40383 \$16 \$11608 \$16 \$153 \$11546 VNB sky130_fd_sc_hd__clkbuf_2
X$40385 \$153 \$11647 \$11452 \$10326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40386 \$153 \$11702 \$11452 \$10467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40388 \$16 \$10467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40390 \$153 \$11454 \$10285 \$11515 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40391 \$16 \$10326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40392 \$16 \$10392 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40394 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$40395 \$153 \$11703 \$11452 \$10446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40396 \$153 \$11610 \$11452 \$10393 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40397 \$153 \$11610 \$10694 \$11515 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40399 \$153 \$11481 \$10560 \$11515 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40401 \$16 \$10446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40402 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$40404 \$16 \$10326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40405 \$153 \$11705 \$11628 \$10393 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40406 \$153 \$11583 \$10466 \$11829 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40407 \$153 \$11584 \$10285 \$11829 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40408 \$153 \$11583 \$11628 \$10326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40411 \$153 \$11361 \$11316 \$10393 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40413 \$153 \$11706 \$11629 \$10393 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40414 \$16 \$11502 \$16 \$153 \$11384 VNB sky130_fd_sc_hd__inv_1
X$40416 \$153 \$11551 \$11316 \$10467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40417 \$16 \$10393 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40419 \$16 \$10467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40420 \$16 \$12612 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40421 \$153 \$11283 \$12612 \$11707 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$40422 \$153 \$11551 \$10587 \$11384 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40423 \$16 \$11502 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40424 \$153 \$11552 \$10376 \$11495 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40426 \$153 \$11677 \$10466 \$11678 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40430 \$16 \$10617 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40431 \$153 \$11708 \$11709 \$10393 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40432 \$153 \$11566 \$11283 \$10617 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40433 \$153 \$11679 \$10466 \$11680 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40434 \$153 \$11566 \$10560 \$11495 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40435 \$16 \$10346 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40438 \$153 \$11710 \$11709 \$10346 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40439 \$16 \$11496 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40440 \$16 \$11585 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40441 \$153 \$11346 \$11585 \$11553 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$40442 \$153 \$11586 \$11681 \$10326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40443 \$153 \$11019 \$10587 \$11516 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40445 \$153 \$11586 \$10466 \$11730 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40446 \$153 \$11711 \$11681 \$10393 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40447 \$16 \$10446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40448 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$40449 \$153 \$10565 \$10815 \$10858 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40451 \$16 \$11627 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40452 \$16 \$10326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40453 \$153 \$11611 \$11587 \$10326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40454 \$16 \$11413 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40456 \$153 \$11106 \$10285 \$11516 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40457 \$16 \$11413 \$16 \$153 \$11731 VNB sky130_fd_sc_hd__inv_1
X$40458 \$16 \$10393 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40459 \$153 \$11020 \$10376 \$11516 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40460 \$153 \$11712 \$11587 \$10393 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40461 \$16 \$11459 \$16 \$153 \$11390 VNB sky130_fd_sc_hd__inv_1
X$40462 \$16 \$11483 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40464 \$153 \$10935 \$10466 \$11516 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40465 \$153 \$11682 \$11587 \$10346 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40466 \$153 \$11152 \$10815 \$11516 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40467 \$153 \$11682 \$10285 \$11731 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40468 \$153 \$11612 \$11588 \$10446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40471 \$16 \$11546 \$11229 \$11556 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$40472 \$16 \$10393 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40474 \$16 \$10346 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40475 \$16 \$10326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40476 \$153 \$11713 \$11588 \$10346 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40477 \$153 \$11589 \$10285 \$11461 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40478 \$153 \$11590 \$10642 \$11461 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40479 \$153 \$11714 \$11648 \$10393 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40481 \$153 \$10424 \$10285 \$10801 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40482 \$153 \$10701 \$10642 \$10801 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40483 \$153 \$11715 \$11648 \$10346 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40484 \$153 \$11023 \$10466 \$11022 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40485 \$16 \$11546 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40487 \$16 \$10617 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40488 \$16 \$10346 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40490 \$153 \$11613 \$11498 \$10617 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40491 \$153 \$11716 \$11498 \$10446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40492 \$153 \$10702 \$10815 \$10741 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40493 \$153 \$10937 \$10560 \$11022 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40495 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$40496 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$40497 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$40498 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$40499 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$40500 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$40501 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$40502 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$40503 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$40504 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$40506 \$16 \$12230 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40507 \$153 \$12939 \$12839 \$12294 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40510 \$153 \$13026 \$13063 \$12158 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40511 \$153 \$12986 \$12412 \$12982 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40512 \$153 \$13026 \$12057 \$12982 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40513 \$153 \$12939 \$12208 \$12828 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40514 \$16 \$12158 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40516 \$16 \$11289 \$12779 \$13027 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$40518 \$153 \$12893 \$12839 \$12236 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40519 \$153 \$13063 \$11432 \$13027 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$40520 \$16 \$12236 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40521 \$153 \$13044 \$12134 \$12982 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40523 \$153 \$12940 \$12839 \$12093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40526 \$16 \$11432 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40527 \$16 \$11289 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40528 \$153 \$13045 \$12229 \$12982 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40529 \$153 \$12987 \$11810 \$12982 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40530 \$16 \$12093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40531 \$153 \$12940 \$12229 \$12828 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40532 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$40533 \$153 \$12988 \$12842 \$12158 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40535 \$16 \$11369 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40537 \$16 \$12003 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40538 \$16 \$11369 \$16 \$153 \$12924 VNB sky130_fd_sc_hd__inv_1
X$40539 \$153 \$12988 \$12057 \$12924 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40540 \$153 \$12910 \$12842 \$12294 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40541 \$153 \$12941 \$12842 \$12152 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40542 \$16 \$11274 \$12779 \$12873 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$40545 \$153 \$12941 \$12209 \$12924 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40546 \$153 \$13046 \$12134 \$12829 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40547 \$153 \$13065 \$12874 \$12152 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40549 \$153 \$12843 \$12874 \$12003 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40550 \$16 \$12152 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40552 \$16 \$12236 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40553 \$16 \$12003 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40555 \$16 \$11274 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40556 \$153 \$12942 \$12874 \$12158 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40557 \$16 \$12013 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40558 \$153 \$13028 \$12874 \$12294 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40559 \$153 \$12942 \$12057 \$12829 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40560 \$16 \$12294 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40561 \$16 \$12230 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40562 \$16 \$12003 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40564 \$16 \$12158 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40566 \$153 \$12989 \$12720 \$12294 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40567 \$153 \$12912 \$12720 \$12003 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40568 \$153 \$13028 \$12208 \$12829 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40569 \$153 \$12989 \$12208 \$12780 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40570 \$153 \$13029 \$12720 \$12230 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40572 \$153 \$12990 \$12209 \$12780 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40573 \$16 \$12003 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40574 \$16 \$11800 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40575 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$40576 \$153 \$13029 \$12412 \$12780 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40577 \$153 \$12925 \$12875 \$12095 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40578 \$16 \$12230 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40579 \$16 \$11897 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40582 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$40583 \$153 \$12943 \$12229 \$12926 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40584 \$16 \$12095 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40585 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$40586 \$153 \$12875 \$11856 \$12927 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$40587 \$153 \$12812 \$11810 \$12926 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40588 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$40589 \$16 \$11856 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40591 \$153 \$12898 \$12057 \$12926 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40593 \$16 \$11240 \$16 \$153 \$12926 VNB sky130_fd_sc_hd__inv_1
X$40594 \$16 \$11240 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40596 \$153 \$12845 \$12921 \$12152 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40597 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$40598 \$153 \$13067 \$12921 \$12003 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40599 \$153 \$12991 \$12921 \$12236 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40600 \$16 \$12152 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40602 \$16 \$12003 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40603 \$153 \$12813 \$12134 \$12579 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40604 \$16 \$11594 \$16 \$153 \$12795 VNB sky130_fd_sc_hd__inv_1
X$40605 \$16 \$12236 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40607 \$153 \$12993 \$10959 \$12992 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$40608 \$16 \$11267 \$12897 \$12945 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$40609 \$153 \$13047 \$12353 \$12795 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40611 \$16 \$10974 \$12897 \$12992 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$40612 \$153 \$12944 \$12208 \$12795 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40614 \$153 \$13068 \$12993 \$12294 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40615 \$16 \$11431 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40616 \$16 \$12152 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40617 \$153 \$12994 \$12708 \$12152 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40618 \$16 \$12294 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40619 \$16 \$12152 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40620 \$16 \$13215 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40622 \$153 \$12946 \$12057 \$12783 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40623 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$40624 \$16 \$11267 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40625 \$153 \$12947 \$12708 \$12230 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40626 \$153 \$12994 \$12209 \$12783 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40627 \$153 \$13160 \$12229 \$13108 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40628 \$16 \$11267 \$16 \$153 \$12783 VNB sky130_fd_sc_hd__inv_1
X$40629 \$16 \$10974 \$16 \$153 \$13108 VNB sky130_fd_sc_hd__inv_1
X$40630 \$153 \$13048 \$12057 \$13215 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40632 \$153 \$12947 \$12412 \$12783 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40633 \$16 \$11432 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40634 \$16 \$12230 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40636 \$16 \$10974 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40637 \$153 \$13030 \$12877 \$12296 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40639 \$153 \$12948 \$12877 \$12259 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40643 \$153 \$13030 \$12359 \$12928 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40644 \$16 \$12259 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40645 \$153 \$12948 \$12307 \$12928 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40646 \$16 \$12296 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40647 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$40648 \$16 \$12295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40649 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$40650 \$153 \$12995 \$12877 \$12101 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40651 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$40653 \$153 \$12995 \$12476 \$12928 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40654 \$16 \$12101 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40655 \$16 \$12241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40656 \$153 \$12901 \$12174 \$12928 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40657 \$16 \$12241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40658 \$153 \$13031 \$12848 \$12241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40660 \$16 \$11369 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40661 \$16 \$11567 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40662 \$16 \$12160 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40663 \$153 \$12949 \$12848 \$12160 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40665 \$16 \$12241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40667 \$16 \$12160 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40668 \$153 \$13031 \$12363 \$12781 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40669 \$153 \$12949 \$12028 \$12781 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40670 \$153 \$13032 \$12848 \$12296 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40672 \$16 \$11274 \$12922 \$12996 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$40674 \$16 \$12083 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40675 \$153 \$12997 \$11190 \$12996 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$40676 \$153 \$13032 \$12359 \$12781 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40677 \$16 \$12296 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40678 \$16 \$11190 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40679 \$16 \$11274 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40680 \$153 \$12929 \$12710 \$12160 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40681 \$16 \$11274 \$16 \$153 \$13071 VNB sky130_fd_sc_hd__inv_1
X$40682 \$16 \$12013 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40683 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$40686 \$153 \$13033 \$12997 \$12083 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40687 \$16 \$12160 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40688 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$40689 \$153 \$12930 \$12710 \$12241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40690 \$153 \$13033 \$12174 \$13071 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40691 \$16 \$12083 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40694 \$153 \$13072 \$12997 \$12295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40695 \$16 \$12241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40697 \$153 \$12950 \$12307 \$12729 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40698 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$40699 \$153 \$12851 \$12765 \$12259 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40700 \$153 \$13034 \$12363 \$13071 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40701 \$16 \$12295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40704 \$16 \$11800 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40705 \$16 \$12259 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40706 \$153 \$12998 \$12765 \$12044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40707 \$16 \$11897 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40708 \$16 \$11800 \$12785 \$13074 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$40709 \$153 \$12998 \$12068 \$12758 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40710 \$153 \$12951 \$12359 \$12758 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40711 \$153 \$13035 \$13042 \$12101 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40713 \$153 \$12852 \$12765 \$12295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40714 \$153 \$12952 \$12174 \$12758 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40715 \$16 \$12083 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40716 \$153 \$13036 \$12307 \$13049 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40717 \$16 \$12295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40718 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$40719 \$153 \$12853 \$12508 \$12044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40720 \$16 \$12101 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40722 \$153 \$13035 \$12476 \$13049 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40723 \$16 \$12160 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40724 \$153 \$12954 \$12307 \$12429 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40725 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$40726 \$16 \$11240 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40727 \$153 \$13075 \$13042 \$12044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40728 \$16 \$12044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40730 \$16 \$11240 \$12785 \$12955 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$40732 \$153 \$12953 \$12155 \$12429 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40733 \$16 \$12044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40734 \$153 \$12816 \$12155 \$12430 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40735 \$153 \$12768 \$12028 \$12430 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40736 \$153 \$13075 \$12068 \$13049 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40738 \$153 \$12999 \$11431 \$12957 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$40739 \$16 \$11240 \$16 \$153 \$13051 VNB sky130_fd_sc_hd__inv_1
X$40742 \$153 \$13050 \$12476 \$13051 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40743 \$16 \$11240 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40744 \$16 \$12160 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40745 \$153 \$13000 \$12879 \$12160 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40746 \$153 \$13076 \$12999 \$12160 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40747 \$16 \$12160 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40751 \$153 \$13000 \$12028 \$12881 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40752 \$153 \$12958 \$12307 \$12881 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40753 \$16 \$11267 \$16 \$153 \$13077 VNB sky130_fd_sc_hd__inv_1
X$40755 \$16 \$12296 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40756 \$153 \$13002 \$12879 \$12083 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40757 \$153 \$12959 \$12155 \$12881 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40758 \$153 \$13001 \$12879 \$12296 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40761 \$153 \$13079 \$12879 \$12044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40762 \$153 \$13001 \$12359 \$12881 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40763 \$16 \$12044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40764 \$153 \$13002 \$12174 \$12881 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40766 \$16 \$12326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40767 \$16 \$12297 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40768 \$153 \$12931 \$12984 \$12326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40771 \$153 \$13003 \$12984 \$12115 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40772 \$153 \$13003 \$12234 \$12932 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40774 \$16 \$12233 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40775 \$153 \$12933 \$12984 \$12233 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40776 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$40777 \$16 \$12219 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40778 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$40780 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$40781 \$153 \$13330 \$11451 \$12960 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$40782 \$16 \$11399 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40783 \$16 \$11399 \$12379 \$12983 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$40784 \$153 \$12984 \$11578 \$12983 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$40785 \$16 \$11399 \$16 \$153 \$12932 VNB sky130_fd_sc_hd__inv_1
X$40787 \$16 \$12298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40788 \$16 \$12326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40789 \$153 \$13037 \$12985 \$12326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40791 \$153 \$12934 \$12985 \$12298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40793 \$153 \$13037 \$12264 \$12935 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40794 \$153 \$13004 \$12736 \$12298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40795 \$16 \$12298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40796 \$16 \$12115 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40798 \$153 \$13083 \$12985 \$12115 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40800 \$153 \$12961 \$12110 \$12787 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40801 \$153 \$13005 \$12217 \$12935 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40802 \$16 \$11824 \$16 \$153 \$12935 VNB sky130_fd_sc_hd__inv_1
X$40804 \$153 \$12985 \$12162 \$13006 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$40805 \$16 \$11824 \$12634 \$13006 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$40807 \$16 \$11824 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40808 \$16 \$11824 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40809 \$16 \$11842 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40810 \$16 \$12219 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40811 \$153 \$12800 \$12309 \$12787 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40812 \$153 \$12857 \$12856 \$12219 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40813 \$16 \$12162 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40814 \$16 \$12009 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40815 \$153 \$13172 \$12309 \$12832 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40816 \$153 \$12962 \$12217 \$12832 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40818 \$153 \$13084 \$12582 \$12832 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40819 \$153 \$12884 \$12603 \$12832 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40820 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$40822 \$153 \$13052 \$12165 \$12832 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40823 \$153 \$12963 \$12264 \$12832 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40824 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$40825 \$16 \$12164 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40826 \$16 \$11214 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40827 \$16 \$12571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40829 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$40830 \$153 \$12859 \$12916 \$12571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40831 \$153 \$13038 \$12264 \$12648 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40832 \$153 \$13173 \$12603 \$12833 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40834 \$16 \$12326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40835 \$153 \$12861 \$12916 \$12326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40836 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$40838 \$16 \$11214 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40840 \$153 \$13053 \$12165 \$12833 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40841 \$153 \$12964 \$12234 \$12833 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40842 \$16 \$12298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40843 \$16 \$12219 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40844 \$16 \$12219 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40845 \$153 \$13007 \$13054 \$12219 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40847 \$153 \$13007 \$12110 \$12648 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40849 \$153 \$13008 \$12670 \$12571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40850 \$153 \$12965 \$12264 \$12671 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40851 \$153 \$13008 \$12309 \$12671 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40852 \$153 \$13009 \$12917 \$12115 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40853 \$16 \$11627 \$12820 \$13086 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$40857 \$153 \$13009 \$12234 \$12863 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40858 \$16 \$12820 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40860 \$16 \$12326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40861 \$153 \$13010 \$12917 \$12326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40862 \$16 \$12297 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40864 \$153 \$13087 \$12917 \$12298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40866 \$16 \$12298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40868 \$153 \$13011 \$12714 \$12298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40869 \$16 \$12298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40871 \$16 \$11798 \$12820 \$13088 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$40872 \$153 \$13011 \$12165 \$12706 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40874 \$16 \$12219 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40876 \$153 \$12936 \$12714 \$12219 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40877 \$153 \$12694 \$12309 \$12706 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40880 \$16 \$12219 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40881 \$153 \$12741 \$12264 \$12706 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40882 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$40883 \$16 \$12571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40884 \$153 \$12834 \$12923 \$12571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40885 \$153 \$13090 \$12923 \$12219 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40887 \$153 \$13091 \$12923 \$12298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40888 \$16 \$12298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40889 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$40890 \$153 \$12774 \$12582 \$12488 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40891 \$16 \$11172 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40892 \$153 \$13090 \$12110 \$12836 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40893 \$16 \$12326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40894 \$153 \$12966 \$12217 \$12836 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40896 \$16 \$12233 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40900 \$153 \$12967 \$12923 \$12326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40901 \$153 \$13039 \$12923 \$12115 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40902 \$153 \$12967 \$12264 \$12836 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40903 \$153 \$13039 \$12234 \$12836 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40904 \$16 \$11385 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40905 \$16 \$12115 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40907 \$16 \$11172 \$16 \$153 \$12836 VNB sky130_fd_sc_hd__inv_1
X$40908 \$16 \$11459 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40911 \$16 \$11172 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40912 \$153 \$13012 \$11578 \$12968 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$40914 \$153 \$13092 \$13012 \$12010 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40915 \$16 \$11578 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40916 \$16 \$11374 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40917 \$16 \$12010 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40918 \$16 \$11399 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40919 \$16 \$12303 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40920 \$16 \$11399 \$16 \$153 \$13093 VNB sky130_fd_sc_hd__inv_1
X$40921 \$153 \$12969 \$13012 \$12303 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40924 \$153 \$12937 \$13012 \$12384 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40925 \$153 \$12969 \$12227 \$13093 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40926 \$16 \$12384 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40927 \$153 \$13094 \$12162 \$13013 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$40928 \$16 \$11824 \$12747 \$13013 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$40930 \$153 \$12837 \$12715 \$11983 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40931 \$16 \$11824 \$16 \$153 \$13056 VNB sky130_fd_sc_hd__inv_1
X$40932 \$16 \$11983 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40933 \$16 \$11824 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40934 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$40935 \$16 \$11842 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40936 \$16 \$11824 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40937 \$153 \$13055 \$11881 \$13056 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40938 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$40939 \$16 \$12351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40940 \$153 \$13014 \$12715 \$12351 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40941 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$40943 \$16 \$11502 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40944 \$153 \$13014 \$12119 \$12824 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40945 \$153 \$12971 \$12179 \$12824 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40946 \$153 \$13057 \$11881 \$13058 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40947 \$16 \$12303 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40948 \$153 \$13095 \$12888 \$12303 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40949 \$16 \$12120 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40951 \$16 \$11983 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40953 \$153 \$12867 \$12888 \$11983 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40954 \$153 \$13040 \$12888 \$12351 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40955 \$153 \$12938 \$12888 \$12384 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40956 \$16 \$12351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40957 \$16 \$12120 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40959 \$153 \$13059 \$12339 \$12838 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40960 \$153 \$12972 \$11942 \$12838 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40961 \$153 \$13096 \$12889 \$12120 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40962 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$40963 \$153 \$13015 \$12119 \$12825 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40965 \$16 \$12287 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40967 \$16 \$11983 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40968 \$16 \$12010 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40970 \$153 \$12973 \$12889 \$11983 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40971 \$153 \$13041 \$12889 \$12287 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40972 \$153 \$12973 \$11881 \$12825 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40973 \$153 \$13060 \$12227 \$12825 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40976 \$153 \$13016 \$12890 \$12351 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40977 \$153 \$13041 \$12339 \$12825 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40978 \$16 \$11496 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40980 \$16 \$11496 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40981 \$16 \$11459 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40983 \$153 \$12679 \$12119 \$12680 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40984 \$153 \$13061 \$12227 \$12907 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40985 \$16 \$11983 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40986 \$153 \$12974 \$11942 \$12907 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40988 \$153 \$13017 \$12890 \$11983 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40989 \$16 \$12120 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$40991 \$153 \$13017 \$11881 \$12907 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40992 \$153 \$12975 \$12179 \$12907 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40993 \$153 \$13099 \$12339 \$12907 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40994 \$153 \$12977 \$12807 \$12303 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40997 \$153 \$13101 \$12807 \$12351 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$40998 \$153 \$12977 \$12227 \$12750 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$40999 \$16 \$12299 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41000 \$153 \$13019 \$12807 \$12299 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41002 \$16 \$11172 \$12678 \$13018 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$41004 \$16 \$12287 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41005 \$16 \$11483 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41006 \$153 \$13019 \$12371 \$12750 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41007 \$153 \$12808 \$11881 \$12750 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41008 \$153 \$13020 \$11280 \$13018 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$41009 \$153 \$12978 \$12339 \$12750 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41010 \$16 \$12287 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41011 \$16 \$12010 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41012 \$153 \$13021 \$12872 \$12287 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41014 \$16 \$12120 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41015 \$153 \$13102 \$13020 \$12120 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41016 \$16 \$11627 \$16 \$153 \$12980 VNB sky130_fd_sc_hd__inv_1
X$41018 \$153 \$13022 \$10694 \$12782 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41019 \$153 \$13103 \$13020 \$12010 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41021 \$153 \$13023 \$12872 \$12010 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41023 \$16 \$12384 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41024 \$16 \$12299 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41026 \$153 \$13043 \$13020 \$12351 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41028 \$153 \$13024 \$12872 \$12384 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41030 \$153 \$13062 \$12339 \$13107 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41031 \$153 \$13025 \$12872 \$12351 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41032 \$153 \$13043 \$12119 \$13107 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41034 \$153 \$11559 \$10587 \$12782 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41035 \$16 \$12351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41036 \$16 \$12782 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41037 \$16 \$11627 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41040 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$41041 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$41042 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$41043 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$41044 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$41045 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$41046 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$41048 \$153 \$12314 \$12208 \$12150 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41050 \$153 \$12304 \$12057 \$12150 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41051 \$153 \$12340 \$12251 \$12152 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41052 \$153 \$12314 \$12251 \$12294 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41054 \$16 \$12152 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41056 \$16 \$12294 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41057 \$153 \$12315 \$12251 \$12230 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41058 \$153 \$12375 \$12353 \$12150 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41059 \$153 \$12304 \$12251 \$12158 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41060 \$16 \$12230 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41061 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$41062 \$16 \$10730 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41064 \$153 \$12151 \$12251 \$12236 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41065 \$16 \$12158 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41066 \$16 \$10764 \$12012 \$12354 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$41067 \$153 \$12355 \$10888 \$12354 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$41068 \$153 \$12091 \$12353 \$12020 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41069 \$16 \$10764 \$16 \$153 \$12386 VNB sky130_fd_sc_hd__inv_1
X$41070 \$16 \$12236 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41071 \$16 \$10888 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41073 \$153 \$12436 \$12251 \$12093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41075 \$153 \$12375 \$12251 \$12095 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41076 \$16 \$10730 \$16 \$153 \$12150 VNB sky130_fd_sc_hd__inv_1
X$41077 \$153 \$12376 \$11810 \$12386 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41078 \$153 \$12305 \$12134 \$12252 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41080 \$153 \$12305 \$12041 \$12236 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41082 \$153 \$12316 \$12041 \$12294 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41083 \$153 \$12316 \$12208 \$12252 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41084 \$153 \$12317 \$12041 \$12152 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41085 \$16 \$10939 \$12012 \$12387 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$41087 \$153 \$12317 \$12209 \$12252 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41088 \$153 \$12318 \$12041 \$12230 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41090 \$153 \$12306 \$11989 \$12294 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41091 \$16 \$12152 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41092 \$16 \$12230 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41093 \$16 \$10939 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41094 \$16 \$10744 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41095 \$16 \$12294 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41099 \$153 \$12388 \$11989 \$12236 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41100 \$153 \$12272 \$11989 \$12230 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41101 \$153 \$12306 \$12208 \$12094 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41102 \$153 \$12253 \$12209 \$12094 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41104 \$16 \$12236 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41105 \$153 \$12273 \$12014 \$12294 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41107 \$153 \$12389 \$12014 \$12230 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41108 \$153 \$12272 \$12412 \$12094 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41109 \$153 \$12388 \$12134 \$12094 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41110 \$16 \$12294 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41111 \$16 \$12230 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41113 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$41115 \$153 \$12341 \$12014 \$12152 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41116 \$153 \$12341 \$12209 \$12004 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41117 \$153 \$12342 \$12096 \$12236 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41118 \$153 \$12255 \$12096 \$12294 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41120 \$153 \$12377 \$12134 \$12578 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41121 \$16 \$12294 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41122 \$16 \$12152 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41123 \$16 \$10413 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41124 \$153 \$12237 \$12096 \$12152 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41125 \$153 \$12390 \$12096 \$12230 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41126 \$16 \$12230 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41127 \$16 \$12152 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41129 \$16 \$12093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41130 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$41131 \$16 \$10825 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41134 \$153 \$12356 \$12172 \$12230 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41135 \$153 \$12274 \$12172 \$12152 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41136 \$16 \$12152 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41137 \$153 \$12274 \$12209 \$12006 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41138 \$16 \$12230 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41139 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$41141 \$153 \$12356 \$12412 \$12006 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41142 \$153 \$12275 \$12172 \$12294 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41143 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$41144 \$16 \$12294 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41145 \$153 \$12391 \$10682 \$12319 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$41146 \$153 \$12275 \$12208 \$12006 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41149 \$153 \$8516 \$12152 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$41150 \$16 \$10732 \$12015 \$12319 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$41151 \$153 \$8670 \$12294 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$41152 \$16 \$8516 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41153 \$16 \$10732 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41154 \$16 \$10732 \$16 \$153 \$12392 VNB sky130_fd_sc_hd__inv_1
X$41155 \$16 \$8670 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41159 \$153 \$8671 \$12230 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$41160 \$153 \$8568 \$12236 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$41161 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41162 \$16 \$10764 \$12159 \$12343 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$41163 \$16 \$8671 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41164 \$16 \$8568 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41165 \$153 \$12357 \$10888 \$12343 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$41166 \$16 \$12134 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41168 \$16 \$10730 \$12159 \$12320 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$41170 \$16 \$10603 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41171 \$16 \$12208 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41174 \$153 \$12276 \$12191 \$12296 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41175 \$153 \$12393 \$12357 \$12295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41177 \$153 \$12276 \$12359 \$12135 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41179 \$153 \$12212 \$12155 \$12135 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41180 \$153 \$12256 \$12307 \$12135 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41181 \$153 \$12393 \$12155 \$12427 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41183 \$153 \$12344 \$12363 \$12135 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41184 \$153 \$12344 \$12191 \$12241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41186 \$16 \$12101 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41187 \$16 \$10764 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41188 \$153 \$12103 \$12476 \$12135 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41190 \$16 \$10730 \$16 \$153 \$12154 VNB sky130_fd_sc_hd__inv_1
X$41191 \$153 \$12173 \$12533 \$12241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41192 \$16 \$12241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41193 \$16 \$10539 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41194 \$16 \$10730 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41196 \$153 \$12239 \$11996 \$12259 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41197 \$16 \$12241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41199 \$153 \$12394 \$11996 \$12241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41200 \$16 \$12259 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41201 \$16 \$12295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41202 \$153 \$12277 \$11996 \$12295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41204 \$153 \$12358 \$11996 \$12296 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41206 \$16 \$12296 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41207 \$153 \$12277 \$12155 \$12238 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41208 \$153 \$12358 \$12359 \$12238 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41209 \$153 \$12321 \$12070 \$12259 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41210 \$16 \$10939 \$12159 \$12395 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$41211 \$153 \$12258 \$12476 \$12104 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41212 \$153 \$12321 \$12307 \$12104 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41214 \$16 \$12259 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41215 \$16 \$11114 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41216 \$16 \$10939 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41219 \$153 \$12231 \$12070 \$12295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41220 \$153 \$12322 \$12070 \$12296 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41221 \$153 \$12322 \$12359 \$12104 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41222 \$16 \$12296 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41225 \$16 \$12241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41227 \$153 \$12323 \$12084 \$12296 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41229 \$153 \$12396 \$12084 \$12295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41230 \$16 \$12296 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41231 \$16 \$12295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41232 \$16 \$10555 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41233 \$16 \$10825 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41235 \$16 \$10825 \$16 \$153 \$12360 VNB sky130_fd_sc_hd__inv_1
X$41237 \$153 \$12278 \$12084 \$12259 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41240 \$153 \$12345 \$12084 \$12241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41241 \$153 \$12278 \$12307 \$12071 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41242 \$153 \$12397 \$12085 \$12241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41243 \$16 \$12259 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41244 \$16 \$12241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41247 \$153 \$12345 \$12363 \$12071 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41248 \$16 \$12241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41249 \$153 \$12361 \$12085 \$12296 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41251 \$16 \$10732 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41252 \$153 \$12279 \$12085 \$12259 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41254 \$16 \$10732 \$12161 \$12260 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$41256 \$153 \$12279 \$12307 \$12007 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41257 \$153 \$12361 \$12359 \$12007 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41258 \$153 \$12240 \$12086 \$12296 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41259 \$153 \$12398 \$12086 \$12295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41260 \$16 \$12295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41261 \$16 \$12296 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41263 \$153 \$12362 \$12308 \$12241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41264 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$41265 \$153 \$12280 \$12086 \$12259 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41267 \$153 \$12362 \$12363 \$12378 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41268 \$153 \$12280 \$12307 \$11869 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41269 \$16 \$10732 \$16 \$153 \$12378 VNB sky130_fd_sc_hd__inv_1
X$41271 \$16 \$12259 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41272 \$16 \$12241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41273 \$16 \$10732 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41274 \$16 \$11594 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41276 \$153 \$12324 \$12308 \$12083 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41277 \$153 \$12242 \$12308 \$12044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41279 \$153 \$12324 \$12174 \$12378 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41280 \$16 \$8416 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41281 \$16 \$12083 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41284 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$41285 \$16 \$12044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41286 \$153 \$8391 \$12241 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$41288 \$153 \$8347 \$12296 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$41289 \$16 \$10383 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41290 \$16 \$8391 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41291 \$16 \$8364 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41293 \$16 \$8347 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41295 \$16 \$8670 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41297 \$153 \$8670 \$12297 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$41298 \$16 \$8671 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41299 \$153 \$8671 \$12571 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$41300 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41301 \$16 \$8516 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41302 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$41305 \$153 \$8516 \$12233 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$41306 \$16 \$11207 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41307 \$16 \$12363 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41308 \$153 \$11698 \$10714 \$11207 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41309 \$153 \$12399 \$12309 \$12690 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41310 \$153 \$8568 \$12298 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$41314 \$16 \$11113 \$12379 \$12364 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$41315 \$153 \$12400 \$11148 \$12364 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$41316 \$16 \$11113 \$16 \$153 \$12325 VNB sky130_fd_sc_hd__inv_1
X$41318 \$16 \$10300 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41319 \$153 \$153 \$12264 \$12243 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41321 \$16 \$10478 \$16 \$153 \$12243 VNB sky130_fd_sc_hd__clkbuf_2
X$41322 \$16 \$12110 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41323 \$153 \$153 \$12603 \$12243 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41325 \$153 \$153 \$12582 \$12243 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41326 \$153 \$153 \$12234 \$12243 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41327 \$153 \$153 \$12309 \$12243 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41328 \$16 \$10478 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41329 \$16 \$12359 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41330 \$16 \$10978 \$12379 \$12401 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$41331 \$16 \$12326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41332 \$153 \$12327 \$12175 \$12326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41333 \$16 \$10978 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41336 \$16 \$11930 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41338 \$16 \$12571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41339 \$153 \$12327 \$12264 \$12216 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41340 \$153 \$12328 \$12175 \$12298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41341 \$153 \$12402 \$12175 \$12571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41342 \$16 \$12298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41344 \$153 \$12262 \$12234 \$12216 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41346 \$153 \$12175 \$10897 \$12380 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$41347 \$16 \$11930 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41348 \$16 \$12297 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41349 \$153 \$12329 \$12175 \$12297 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41350 \$16 \$11013 \$12379 \$12403 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$41351 \$16 \$10739 \$12379 \$12380 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$41353 \$153 \$12329 \$12582 \$12216 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41354 \$153 \$12244 \$12175 \$12233 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41355 \$16 \$12326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41356 \$153 \$12365 \$12163 \$12326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41357 \$16 \$12233 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41358 \$153 \$12310 \$12309 \$12156 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41361 \$153 \$12263 \$12110 \$12156 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41362 \$153 \$12281 \$12163 \$12298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41363 \$153 \$12365 \$12264 \$12156 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41365 \$153 \$12330 \$12163 \$12297 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41367 \$153 \$12331 \$12603 \$12156 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41369 \$153 \$12330 \$12582 \$12156 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41370 \$153 \$12331 \$12163 \$12233 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41371 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$41372 \$16 \$12164 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41373 \$153 \$12346 \$12113 \$12164 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41375 \$16 \$12115 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41376 \$16 \$12298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41377 \$16 \$12326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41379 \$153 \$12282 \$12113 \$12326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41380 \$153 \$12366 \$12113 \$12298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41381 \$153 \$12283 \$12075 \$12164 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41382 \$153 \$12366 \$12165 \$12200 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41386 \$153 \$12141 \$12110 \$11999 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41387 \$153 \$12455 \$12075 \$12233 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41388 \$153 \$12177 \$12245 \$12332 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$41389 \$16 \$10597 \$12166 \$12332 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$41391 \$153 \$12367 \$12177 \$12233 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41392 \$16 \$12164 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41394 \$153 \$12284 \$12177 \$12164 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41395 \$153 \$12367 \$12603 \$12117 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41396 \$153 \$12284 \$12217 \$12117 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41397 \$16 \$10597 \$16 \$153 \$12117 VNB sky130_fd_sc_hd__inv_1
X$41398 \$16 \$12245 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41399 \$16 \$10597 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41400 \$16 \$12571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41401 \$16 \$12297 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41404 \$153 \$12285 \$12118 \$12297 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41405 \$153 \$12368 \$12118 \$12571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41408 \$153 \$12285 \$12582 \$12246 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41409 \$153 \$12368 \$12309 \$12246 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41413 \$16 \$12233 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41414 \$16 \$12326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41415 \$153 \$12286 \$12118 \$12233 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41416 \$153 \$12369 \$12118 \$12326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41417 \$153 \$12286 \$12603 \$12246 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41418 \$153 \$12369 \$12264 \$12246 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41419 \$16 \$10853 \$16 \$153 \$12333 VNB sky130_fd_sc_hd__inv_1
X$41422 \$16 \$12348 \$11747 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$41423 \$153 \$10383 \$12287 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$41424 \$153 \$12381 \$12603 \$12333 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41425 \$16 \$10978 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41426 \$16 \$12167 \$10615 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$41428 \$16 \$12168 \$16 \$153 \$12348 VNB sky130_fd_sc_hd__clkbuf_2
X$41429 \$16 \$8340 \$16 \$153 \$12168 VNB sky130_fd_sc_hd__clkbuf_2
X$41430 \$16 \$10478 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41431 \$16 \$10478 \$16 \$153 \$12405 VNB sky130_fd_sc_hd__clkbuf_2
X$41432 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41434 \$16 \$8347 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41435 \$16 \$12168 \$16 \$153 \$12311 VNB sky130_fd_sc_hd__clkbuf_2
X$41436 \$16 \$12311 \$12347 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$41438 \$16 \$12311 \$11148 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$41439 \$16 \$12311 \$11578 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$41440 \$153 \$8347 \$12303 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$41441 \$16 \$12311 \$11451 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$41442 \$16 \$12311 \$12406 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$41443 \$16 \$12311 \$11015 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$41444 \$16 \$12311 \$10897 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$41445 \$16 \$12311 \$10780 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$41446 \$16 \$10978 \$12459 \$12407 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$41447 \$153 \$8391 \$12351 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$41449 \$16 \$8391 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41451 \$153 \$12178 \$11148 \$12334 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$41453 \$153 \$12370 \$12178 \$12303 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41454 \$16 \$11113 \$12459 \$12334 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$41455 \$16 \$11113 \$16 \$153 \$12247 VNB sky130_fd_sc_hd__inv_1
X$41457 \$153 \$12248 \$12178 \$12287 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41458 \$153 \$12370 \$12227 \$12247 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41459 \$153 \$12382 \$12227 \$12423 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41461 \$16 \$12299 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41462 \$153 \$12335 \$12178 \$12299 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41463 \$16 \$11013 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41464 \$16 \$12347 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41466 \$16 \$12351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41467 \$153 \$12335 \$12371 \$12247 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41468 \$153 \$12288 \$12178 \$12351 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41469 \$153 \$12170 \$10897 \$12336 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$41470 \$16 \$10739 \$12459 \$12336 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$41471 \$153 \$12300 \$12170 \$12303 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41473 \$153 \$12249 \$12170 \$12299 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41474 \$153 \$12383 \$12119 \$12337 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41475 \$16 \$11013 \$16 \$153 \$12337 VNB sky130_fd_sc_hd__inv_1
X$41476 \$16 \$12299 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41477 \$153 \$12289 \$12170 \$12384 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41478 \$16 \$11013 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41479 \$16 \$10897 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41480 \$16 \$12287 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41482 \$153 \$12301 \$12170 \$12287 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41483 \$153 \$12300 \$12227 \$12121 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41484 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$41485 \$153 \$12289 \$12179 \$12121 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41486 \$16 \$12287 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41487 \$16 \$12303 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41488 \$153 \$12372 \$12087 \$12287 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41491 \$153 \$12338 \$12087 \$12303 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41492 \$153 \$12349 \$12087 \$12384 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41493 \$153 \$12301 \$12339 \$12121 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41494 \$153 \$12312 \$12180 \$12303 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41496 \$153 \$12338 \$12227 \$12147 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41497 \$16 \$10736 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41498 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$41499 \$153 \$12312 \$12227 \$12302 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41500 \$16 \$12120 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41501 \$153 \$12350 \$12180 \$12120 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41502 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$41505 \$16 \$11983 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41506 \$153 \$12350 \$12182 \$12302 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41507 \$153 \$12267 \$11942 \$12302 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41509 \$16 \$12384 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41510 \$153 \$12126 \$11942 \$12147 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41511 \$153 \$12290 \$12088 \$12384 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41512 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$41516 \$16 \$12287 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41517 \$153 \$12291 \$12088 \$12120 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41519 \$153 \$12408 \$12227 \$12127 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41521 \$153 \$12409 \$12245 \$12313 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$41522 \$16 \$10597 \$12018 \$12313 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$41524 \$16 \$10597 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41526 \$153 \$12291 \$12182 \$12127 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41527 \$16 \$12351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41528 \$153 \$12269 \$12179 \$11958 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41529 \$16 \$10597 \$16 \$153 \$12521 VNB sky130_fd_sc_hd__inv_1
X$41530 \$16 \$10853 \$16 \$153 \$11958 VNB sky130_fd_sc_hd__inv_1
X$41531 \$153 \$12374 \$12089 \$12351 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41533 \$153 \$12292 \$12089 \$12303 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41535 \$153 \$12373 \$10960 \$12410 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$41536 \$153 \$12038 \$12089 \$12287 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41538 \$16 \$12010 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41539 \$153 \$12352 \$12373 \$12010 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41540 \$16 \$11776 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41541 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$41543 \$16 \$12287 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41544 \$16 \$12303 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41545 \$153 \$12271 \$12339 \$12011 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41546 \$153 \$12374 \$12119 \$11958 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41548 \$153 \$12493 \$11881 \$12411 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41549 \$153 \$12293 \$12037 \$12303 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41550 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$41553 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$41554 \$153 \$12293 \$12227 \$12011 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41555 \$153 \$12385 \$12227 \$12411 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41556 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$41557 \$153 \$11928 \$10560 \$11926 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41558 \$153 \$11715 \$10285 \$11926 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41559 \$153 \$11793 \$10376 \$11926 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41560 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$41563 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$41564 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$41565 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$41566 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$41567 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$41568 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$41569 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$41571 \$16 \$12152 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41572 \$153 \$12809 \$12839 \$12152 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41574 \$153 \$12809 \$12209 \$12828 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41575 \$153 \$12790 \$12209 \$12512 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41577 \$16 \$12158 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41579 \$153 \$12839 \$11720 \$12791 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$41580 \$16 \$11720 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41581 \$153 \$12840 \$12839 \$12003 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41582 \$153 \$12841 \$12353 \$12828 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41583 \$153 \$12840 \$11810 \$12828 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41584 \$16 \$12236 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41586 \$153 \$12810 \$12842 \$12236 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41587 \$153 \$12842 \$11567 \$12792 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$41588 \$16 \$12230 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41589 \$153 \$12874 \$11190 \$12873 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$41591 \$153 \$12843 \$11810 \$12829 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41593 \$153 \$12894 \$12353 \$12829 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41594 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$41596 \$153 \$12844 \$12412 \$12829 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41597 \$16 \$11274 \$16 \$153 \$12829 VNB sky130_fd_sc_hd__inv_1
X$41598 \$16 \$12093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41599 \$16 \$11274 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41600 \$153 \$12811 \$12720 \$12093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41601 \$153 \$12811 \$12229 \$12780 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41604 \$16 \$12093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41605 \$16 \$11297 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41607 \$153 \$12794 \$12353 \$12780 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41608 \$153 \$12812 \$12875 \$12003 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41609 \$16 \$12003 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41611 \$153 \$12722 \$12209 \$12413 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41612 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$41613 \$153 \$12845 \$12209 \$12795 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41615 \$153 \$12659 \$12134 \$12413 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41616 \$16 \$11240 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41618 \$153 \$12813 \$12514 \$12236 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41619 \$16 \$12236 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41620 \$153 \$12796 \$12412 \$12579 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41622 \$16 \$11594 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41623 \$153 \$12591 \$11810 \$12579 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41624 \$16 \$11689 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41627 \$16 \$10959 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41628 \$16 \$12230 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41629 \$153 \$12846 \$12708 \$12294 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41630 \$16 \$12294 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41631 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$41632 \$153 \$12725 \$12209 \$12392 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41633 \$153 \$12846 \$12208 \$12783 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41634 \$153 \$12797 \$11810 \$12783 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41636 \$16 \$11720 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41638 \$153 \$12877 \$11720 \$12876 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$41639 \$16 \$11636 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41640 \$16 \$12044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41641 \$153 \$12814 \$12877 \$12295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41642 \$16 \$12259 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41643 \$16 \$12295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41644 \$16 \$12295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41645 \$153 \$12815 \$12615 \$12241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41647 \$16 \$12241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41649 \$16 \$12083 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41650 \$153 \$12815 \$12363 \$12641 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41651 \$153 \$12847 \$12028 \$12928 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41653 \$153 \$12784 \$12848 \$12101 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41654 \$153 \$12878 \$12848 \$12044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41657 \$153 \$12849 \$12174 \$12781 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41658 \$153 \$12594 \$12155 \$12154 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41659 \$16 \$12581 \$16 \$153 \$12922 VNB sky130_fd_sc_hd__clkbuf_2
X$41660 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$41661 \$153 \$12850 \$12155 \$12729 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41663 \$153 \$12764 \$12359 \$12498 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41664 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$41666 \$16 \$11364 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41668 \$153 \$12830 \$12359 \$12729 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41669 \$16 \$12259 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41670 \$16 \$12296 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41671 \$153 \$12645 \$12765 \$12101 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41672 \$153 \$12851 \$12307 \$12758 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41673 \$153 \$12766 \$12028 \$12758 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41674 \$16 \$12101 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41675 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$41677 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$41678 \$153 \$12852 \$12155 \$12758 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41679 \$153 \$12703 \$12508 \$12101 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41680 \$16 \$12101 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41681 \$16 \$12295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41682 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$41683 \$153 \$12853 \$12068 \$12429 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41684 \$16 \$11689 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41685 \$16 \$10974 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41686 \$16 \$10959 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41687 \$16 \$11267 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41689 \$153 \$12816 \$12502 \$12295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41690 \$16 \$12160 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41691 \$16 \$12295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41692 \$153 \$12621 \$10959 \$12831 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$41693 \$16 \$10974 \$12785 \$12831 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$41695 \$153 \$12880 \$12879 \$12101 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41697 \$153 \$12665 \$12028 \$12704 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41698 \$16 \$11594 \$16 \$153 \$12881 VNB sky130_fd_sc_hd__inv_1
X$41699 \$16 \$12101 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41701 \$16 \$12083 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41702 \$153 \$12817 \$12621 \$12083 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41703 \$153 \$12817 \$12174 \$12704 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41704 \$153 \$12596 \$12363 \$12704 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41705 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$41706 \$16 \$12326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41708 \$153 \$12882 \$12711 \$12326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41709 \$153 \$12854 \$12234 \$12690 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41711 \$16 \$12219 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41712 \$16 \$12298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41713 \$153 \$12818 \$12711 \$12298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41714 \$153 \$12855 \$12110 \$12690 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41716 \$153 \$12819 \$12736 \$12297 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41717 \$153 \$12818 \$12165 \$12690 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41718 \$153 \$12819 \$12582 \$12787 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41720 \$153 \$12883 \$12736 \$12164 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41721 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$41725 \$16 \$10854 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41726 \$16 \$12233 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41727 \$153 \$12884 \$12856 \$12233 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41728 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$41729 \$153 \$12857 \$12110 \$12832 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41730 \$16 \$11502 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41732 \$153 \$12856 \$11604 \$12858 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$41733 \$16 \$11502 \$12634 \$12858 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$41736 \$153 \$12916 \$11216 \$12885 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$41737 \$153 \$12859 \$12309 \$12833 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41739 \$153 \$12860 \$12309 \$12648 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41740 \$153 \$12737 \$12603 \$12432 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41741 \$153 \$12861 \$12264 \$12833 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41742 \$16 \$12600 \$16 \$153 \$12820 VNB sky130_fd_sc_hd__clkbuf_2
X$41745 \$16 \$12571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41747 \$153 \$12669 \$12217 \$12671 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41748 \$153 \$12862 \$12110 \$12671 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41750 \$16 \$11627 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41751 \$153 \$12917 \$11585 \$12886 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$41752 \$153 \$12739 \$12603 \$12671 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41753 \$153 \$12864 \$12217 \$12863 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41756 \$16 \$12820 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41757 \$153 \$12627 \$12217 \$12706 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41758 \$16 \$11413 \$12820 \$12801 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$41760 \$153 \$12821 \$12714 \$12297 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41761 \$153 \$12821 \$12582 \$12706 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41762 \$16 \$12219 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41763 \$16 \$11413 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41764 \$153 \$12673 \$12309 \$12488 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41766 \$16 \$12297 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41768 \$153 \$12802 \$12110 \$12488 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41769 \$16 \$10409 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41771 \$16 \$12820 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41772 \$16 \$12326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41773 \$153 \$12923 \$11280 \$12887 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$41774 \$153 \$12835 \$12582 \$12836 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41775 \$153 \$12834 \$12309 \$12836 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41776 \$16 \$11280 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41777 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$41780 \$16 \$11983 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41782 \$153 \$12776 \$12675 \$12010 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41783 \$153 \$12803 \$12371 \$12650 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41784 \$16 \$12010 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41785 \$153 \$12822 \$12675 \$12384 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41786 \$153 \$12822 \$12179 \$12650 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41788 \$16 \$12384 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41789 \$153 \$12823 \$12715 \$12120 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41790 \$153 \$12823 \$12182 \$12824 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41791 \$153 \$12837 \$11881 \$12824 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41792 \$16 \$10831 \$16 \$153 \$12824 VNB sky130_fd_sc_hd__inv_1
X$41793 \$153 \$12888 \$11604 \$12865 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$41795 \$16 \$11502 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41797 \$16 \$12351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41799 \$16 \$12010 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41800 \$16 \$11502 \$16 \$153 \$12838 VNB sky130_fd_sc_hd__inv_1
X$41801 \$153 \$12866 \$12182 \$12838 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41802 \$153 \$12867 \$11881 \$12838 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41804 \$16 \$11216 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41805 \$16 \$11214 \$12747 \$12868 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$41806 \$153 \$12889 \$11216 \$12868 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$41807 \$16 \$11214 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41808 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$41809 \$16 \$11214 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41811 \$153 \$12869 \$12179 \$12825 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41812 \$16 \$11214 \$16 \$153 \$12825 VNB sky130_fd_sc_hd__inv_1
X$41813 \$153 \$12372 \$12339 \$12147 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41815 \$16 \$11585 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41816 \$153 \$12890 \$11585 \$12870 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$41817 \$16 \$11496 \$12678 \$12870 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$41818 \$16 \$11413 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41819 \$153 \$12804 \$12339 \$12680 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41820 \$16 \$12384 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41823 \$16 \$11413 \$12678 \$12806 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$41824 \$153 \$12805 \$12227 \$12680 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41825 \$153 \$12788 \$12635 \$12010 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41826 \$153 \$12826 \$12807 \$12384 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41827 \$153 \$12826 \$12179 \$12750 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41829 \$153 \$12871 \$12807 \$12120 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41830 \$153 \$12871 \$12182 \$12750 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41831 \$16 \$11983 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41832 \$153 \$12762 \$12872 \$11983 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41833 \$153 \$11173 \$10587 \$11322 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41834 \$16 \$12120 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41835 \$16 \$12010 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41837 \$153 \$11135 \$10466 \$11322 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41838 \$153 \$12752 \$12182 \$12654 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41839 \$153 \$12789 \$12636 \$12351 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41840 \$153 \$12827 \$12872 \$12303 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41841 \$16 \$12782 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41842 \$16 \$12782 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41845 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$41846 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$41847 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$41848 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$41850 \$153 \$12891 \$12839 \$12230 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41853 \$153 \$12891 \$12412 \$12828 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41854 \$153 \$12892 \$12839 \$12158 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41855 \$153 \$12892 \$12057 \$12828 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41856 \$16 \$11636 \$16 \$153 \$12828 VNB sky130_fd_sc_hd__inv_1
X$41857 \$153 \$12893 \$12134 \$12828 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41858 \$16 \$11636 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41859 \$16 \$11636 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41860 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$41863 \$153 \$12841 \$12839 \$12095 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41864 \$16 \$12003 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41865 \$16 \$12095 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41866 \$153 \$12911 \$12842 \$12003 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41867 \$153 \$12910 \$12208 \$12924 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41868 \$153 \$12911 \$11810 \$12924 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41869 \$16 \$12294 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41871 \$153 \$12810 \$12134 \$12924 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41872 \$16 \$12152 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41873 \$153 \$12894 \$12874 \$12095 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41874 \$16 \$12095 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41876 \$153 \$12895 \$12874 \$12093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41877 \$153 \$12895 \$12229 \$12829 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41880 \$153 \$12896 \$12720 \$12158 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41881 \$153 \$12896 \$12057 \$12780 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41882 \$153 \$12912 \$11810 \$12780 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41883 \$16 \$12564 \$16 \$153 \$12897 VNB sky130_fd_sc_hd__clkbuf_2
X$41885 \$153 \$12943 \$12875 \$12093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41887 \$16 \$12093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41889 \$153 \$12925 \$12353 \$12926 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41890 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$41891 \$153 \$12898 \$12875 \$12158 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41892 \$16 \$11240 \$12897 \$12927 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$41893 \$16 \$12158 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41894 \$153 \$12944 \$12921 \$12294 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41895 \$16 \$12294 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41898 \$153 \$12921 \$11689 \$12913 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$41899 \$153 \$12708 \$11431 \$12945 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$41900 \$16 \$12158 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41901 \$153 \$12946 \$12708 \$12158 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41902 \$153 \$12660 \$12134 \$12392 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41904 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$41905 \$16 \$12095 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41906 \$153 \$12899 \$12708 \$12095 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41907 \$153 \$12899 \$12353 \$12783 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41908 \$16 \$11636 \$12922 \$12876 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$41909 \$16 \$11636 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41910 \$153 \$12900 \$12877 \$12044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41911 \$16 \$11636 \$16 \$153 \$12928 VNB sky130_fd_sc_hd__inv_1
X$41913 \$153 \$12900 \$12068 \$12928 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41914 \$153 \$12814 \$12155 \$12928 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41916 \$153 \$12901 \$12877 \$12083 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41917 \$153 \$12847 \$12877 \$12160 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41918 \$16 \$11369 \$12922 \$12914 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$41920 \$153 \$12848 \$11567 \$12914 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$41921 \$153 \$12849 \$12848 \$12083 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41922 \$153 \$12878 \$12068 \$12781 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41924 \$153 \$12850 \$12710 \$12295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41926 \$153 \$12929 \$12028 \$12729 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41927 \$16 \$12295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41928 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$41929 \$153 \$12950 \$12710 \$12259 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41930 \$153 \$12830 \$12710 \$12296 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41931 \$153 \$12930 \$12363 \$12729 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41933 \$153 \$12951 \$12765 \$12296 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41934 \$16 \$12296 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41935 \$16 \$12044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41936 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$41937 \$153 \$12952 \$12765 \$12083 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41939 \$153 \$12953 \$12508 \$12295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41941 \$153 \$12954 \$12508 \$12259 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41942 \$16 \$12259 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41944 \$16 \$11856 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41945 \$153 \$12956 \$11856 \$12955 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$41946 \$16 \$11431 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41947 \$16 \$11267 \$12785 \$12957 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$41948 \$153 \$12879 \$11689 \$12915 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$41950 \$153 \$12734 \$12363 \$12430 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41951 \$153 \$12958 \$12879 \$12259 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41952 \$16 \$12259 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41953 \$153 \$12880 \$12476 \$12881 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41954 \$153 \$12959 \$12879 \$12295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41955 \$16 \$12295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41956 \$16 \$12241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41958 \$153 \$12770 \$12879 \$12241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41959 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$41960 \$16 \$12115 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41961 \$16 \$12115 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41962 \$153 \$12854 \$12711 \$12115 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41963 \$153 \$12931 \$12264 \$12932 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41964 \$16 \$11374 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41965 \$16 \$11374 \$12379 \$12960 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$41967 \$153 \$12855 \$12711 \$12219 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41968 \$153 \$12933 \$12603 \$12932 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41970 \$16 \$12233 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41971 \$153 \$12786 \$12736 \$12233 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41972 \$153 \$12934 \$12165 \$12935 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41973 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$41975 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$41977 \$16 \$12219 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41978 \$153 \$12961 \$12736 \$12219 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41979 \$153 \$12883 \$12217 \$12787 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41981 \$16 \$12164 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41982 \$153 \$12962 \$12856 \$12164 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41984 \$16 \$12326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41986 \$16 \$11502 \$16 \$153 \$12832 VNB sky130_fd_sc_hd__inv_1
X$41987 \$153 \$12963 \$12856 \$12326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41989 \$16 \$11214 \$12634 \$12885 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$41990 \$153 \$12902 \$12916 \$12164 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41991 \$153 \$12902 \$12217 \$12833 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$41993 \$16 \$12115 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$41994 \$16 \$11214 \$16 \$153 \$12833 VNB sky130_fd_sc_hd__inv_1
X$41996 \$153 \$12964 \$12916 \$12115 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41997 \$153 \$12862 \$12670 \$12219 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41998 \$153 \$12965 \$12670 \$12326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$41999 \$16 \$12326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42000 \$16 \$12115 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42001 \$16 \$12820 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42002 \$16 \$12164 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42004 \$16 \$11496 \$12820 \$12886 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$42005 \$16 \$11496 \$16 \$153 \$12863 VNB sky130_fd_sc_hd__inv_1
X$42006 \$153 \$12864 \$12917 \$12164 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42007 \$16 \$11496 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42009 \$16 \$12233 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42010 \$153 \$12903 \$12714 \$12233 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42011 \$153 \$12903 \$12603 \$12706 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42012 \$16 \$11413 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42015 \$16 \$12297 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42016 \$153 \$12936 \$12110 \$12706 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42018 \$153 \$12835 \$12923 \$12297 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42019 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$42020 \$16 \$12164 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42021 \$153 \$12966 \$12923 \$12164 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42022 \$16 \$11172 \$12820 \$12887 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$42026 \$153 \$12904 \$12923 \$12233 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42027 \$153 \$12904 \$12603 \$12836 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42028 \$16 \$11399 \$12459 \$12968 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$42029 \$153 \$12918 \$11451 \$12919 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$42030 \$16 \$11374 \$12459 \$12919 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$42031 \$16 \$11399 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42032 \$16 \$11451 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42033 \$16 \$12120 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42036 \$153 \$12970 \$12675 \$12120 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42037 \$153 \$12937 \$12179 \$13093 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42038 \$16 \$12299 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42039 \$153 \$12905 \$12715 \$12299 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42040 \$153 \$12905 \$12371 \$12824 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42042 \$16 \$12384 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42044 \$153 \$12971 \$12715 \$12384 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42045 \$16 \$11502 \$12747 \$12865 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$42046 \$153 \$12866 \$12888 \$12120 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42048 \$16 \$12384 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42049 \$153 \$12972 \$12888 \$12010 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42052 \$153 \$12938 \$12179 \$12838 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42053 \$16 \$12384 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42054 \$153 \$12869 \$12889 \$12384 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42055 \$153 \$12906 \$12889 \$12010 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42056 \$153 \$12906 \$11942 \$12825 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42058 \$16 \$12351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42061 \$16 \$12010 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42062 \$153 \$12974 \$12890 \$12010 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42063 \$16 \$11496 \$16 \$153 \$12907 VNB sky130_fd_sc_hd__inv_1
X$42065 \$153 \$12975 \$12890 \$12384 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42066 \$16 \$12010 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42067 \$16 \$11459 \$12678 \$12976 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$42069 \$153 \$12920 \$11942 \$12750 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42071 \$153 \$12920 \$12807 \$12010 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42072 \$16 \$12010 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42073 \$153 \$12978 \$12807 \$12287 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42074 \$16 \$11798 \$12678 \$12979 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$42075 \$16 \$11921 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42076 \$153 \$12872 \$11776 \$12908 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$42079 \$153 \$11153 \$10376 \$11322 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42080 \$16 \$11627 \$12678 \$12908 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$42081 \$153 \$12909 \$12872 \$12120 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42082 \$153 \$12683 \$11881 \$12654 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42083 \$153 \$12981 \$12872 \$12299 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42086 \$153 \$11462 \$10642 \$12782 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42087 \$153 \$11558 \$10285 \$12782 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42089 \$153 \$11716 \$10376 \$12782 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42090 \$16 \$12782 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42091 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$42092 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$42093 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$42094 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$42095 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$42096 \$16 \$12152 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42097 \$153 \$13212 \$13063 \$12152 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42098 \$153 \$13295 \$13213 \$12158 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42100 \$153 \$13212 \$12209 \$12982 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42102 \$153 \$13266 \$13213 \$12093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42104 \$153 \$13214 \$13130 \$12003 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42105 \$153 \$13214 \$11810 \$13239 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42106 \$16 \$12003 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42107 \$16 \$12093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42109 \$153 \$13267 \$13130 \$12093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42111 \$153 \$13268 \$13250 \$12093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42112 \$153 \$13296 \$13250 \$12158 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42113 \$16 \$11794 \$12779 \$13192 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$42114 \$16 \$12158 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42116 \$153 \$13065 \$12209 \$12829 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42117 \$16 \$12093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42118 \$153 \$13269 \$13115 \$12158 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42119 \$16 \$12158 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42121 \$153 \$13193 \$12229 \$13194 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42123 \$153 \$13270 \$13188 \$12158 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42125 \$153 \$13157 \$12134 \$12780 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42126 \$153 \$13195 \$12229 \$13216 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42128 \$153 \$13271 \$12875 \$12236 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42129 \$153 \$13272 \$11637 \$13251 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$42130 \$16 \$11485 \$12897 \$13251 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$42131 \$16 \$12236 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42133 \$153 \$13217 \$13272 \$12003 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42134 \$153 \$13217 \$11810 \$13343 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42135 \$153 \$13133 \$12229 \$12795 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42137 \$153 \$13305 \$12190 \$13297 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$42138 \$16 \$11795 \$12897 \$13273 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$42139 \$16 \$12158 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42141 \$16 \$11795 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42142 \$16 \$12190 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42143 \$153 \$13306 \$12993 \$12003 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42144 \$153 \$13159 \$12057 \$13108 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42145 \$16 \$12003 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42147 \$153 \$13218 \$12993 \$12230 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42148 \$16 \$12230 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42150 \$16 \$11898 \$12922 \$13274 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$42152 \$153 \$13218 \$12412 \$13108 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42153 \$16 \$11289 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42154 \$16 \$11898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42155 \$153 \$13219 \$13118 \$12259 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42157 \$153 \$13219 \$12307 \$13105 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42158 \$153 \$13459 \$12208 \$13215 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42159 \$16 \$13215 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42161 \$16 \$11987 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42162 \$16 \$12083 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42164 \$153 \$13252 \$12028 \$13105 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42165 \$153 \$13220 \$11987 \$13221 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$42166 \$153 \$13196 \$13220 \$12083 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42167 \$153 \$13374 \$12359 \$13222 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42169 \$16 \$11794 \$12922 \$13253 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$42170 \$16 \$12083 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42172 \$153 \$13275 \$11888 \$13253 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$42173 \$153 \$13276 \$12013 \$13189 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$42174 \$153 \$13163 \$12028 \$13071 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42176 \$153 \$13254 \$12476 \$13327 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42177 \$153 \$13277 \$12476 \$13240 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42179 \$153 \$13034 \$12997 \$12241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42180 \$153 \$13299 \$12359 \$13240 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42181 \$16 \$12241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42183 \$16 \$12083 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42184 \$16 \$11485 \$12785 \$13197 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$42186 \$153 \$13223 \$13190 \$12083 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42187 \$16 \$12083 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42188 \$16 \$11800 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42190 \$153 \$13223 \$12174 \$13241 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42191 \$153 \$13278 \$12068 \$13241 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42192 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$42193 \$16 \$11995 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42194 \$153 \$13224 \$11995 \$13255 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$42195 \$153 \$13279 \$12174 \$13242 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42196 \$153 \$13166 \$12155 \$13049 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42199 \$153 \$13256 \$12476 \$13242 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42200 \$153 \$13280 \$12956 \$12296 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42201 \$153 \$13300 \$12956 \$12044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42202 \$153 \$13281 \$12028 \$13051 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42203 \$16 \$12044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42205 \$16 \$11814 \$16 \$153 \$13243 VNB sky130_fd_sc_hd__inv_1
X$42207 \$16 \$12101 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42208 \$153 \$13282 \$12999 \$12295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42209 \$153 \$13225 \$12999 \$12296 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42210 \$153 \$13225 \$12359 \$13077 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42211 \$153 \$13257 \$12363 \$13243 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42213 \$16 \$12571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42215 \$153 \$13198 \$12984 \$12571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42216 \$153 \$13283 \$12264 \$13244 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42218 \$153 \$13199 \$12165 \$12932 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42219 \$153 \$13226 \$13258 \$12219 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42220 \$16 \$12219 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42222 \$16 \$12571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42225 \$16 \$12219 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42226 \$153 \$13227 \$12985 \$12571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42227 \$153 \$13227 \$12309 \$12935 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42228 \$153 \$13004 \$12165 \$12787 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42229 \$153 \$13201 \$12582 \$12935 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42231 \$153 \$13301 \$12110 \$13245 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42233 \$153 \$13315 \$12009 \$13259 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$42234 \$16 \$11772 \$12634 \$13259 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$42236 \$153 \$13284 \$13316 \$12115 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42237 \$16 \$12298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42238 \$16 \$12219 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42239 \$153 \$13317 \$13316 \$12219 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42241 \$16 \$12032 \$16 \$153 \$13302 VNB sky130_fd_sc_hd__inv_1
X$42242 \$153 \$13285 \$12169 \$13228 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$42243 \$16 \$12032 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42244 \$16 \$12169 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42246 \$16 \$12219 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42247 \$153 \$13229 \$13285 \$12219 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42248 \$153 \$13229 \$12110 \$13203 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42249 \$16 \$12115 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42250 \$16 \$11627 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42251 \$16 \$12298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42253 \$153 \$12626 \$13054 \$12298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42255 \$153 \$13146 \$12582 \$12863 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42256 \$153 \$13287 \$13260 \$12219 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42257 \$153 \$13286 \$12217 \$13109 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42258 \$16 \$12326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42259 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$42262 \$16 \$11798 \$16 \$153 \$13109 VNB sky130_fd_sc_hd__inv_1
X$42263 \$16 \$11798 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42264 \$16 \$12326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42265 \$153 \$13231 \$13110 \$12326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42267 \$153 \$13231 \$12264 \$13205 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42268 \$153 \$13087 \$12165 \$12863 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42269 \$16 \$12219 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42270 \$16 \$11483 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42271 \$153 \$13261 \$12165 \$13232 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42273 \$16 \$12820 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42274 \$153 \$13176 \$12110 \$13149 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42275 \$153 \$13288 \$12582 \$13149 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42276 \$16 \$11459 \$12820 \$13122 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$42278 \$16 \$12233 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42279 \$153 \$13233 \$13175 \$12233 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42280 \$153 \$13233 \$12603 \$13149 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42281 \$16 \$11546 \$16 \$153 \$13232 VNB sky130_fd_sc_hd__inv_1
X$42284 \$153 \$13234 \$13012 \$12287 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42285 \$153 \$13234 \$12339 \$13093 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42287 \$16 \$12120 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42288 \$153 \$13235 \$13012 \$12351 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42289 \$153 \$13235 \$12119 \$13093 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42290 \$16 \$12384 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42292 \$153 \$13320 \$13094 \$12384 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42294 \$16 \$11930 \$12747 \$13124 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$42295 \$16 \$11983 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42296 \$153 \$13057 \$13152 \$11983 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42297 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$42298 \$16 \$11772 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42299 \$153 \$13303 \$12179 \$13058 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42300 \$16 \$12120 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42302 \$153 \$13236 \$13180 \$12120 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42303 \$153 \$13236 \$12182 \$13181 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42304 \$153 \$13262 \$12119 \$13181 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42305 \$153 \$13289 \$12198 \$13246 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$42306 \$16 \$12032 \$12747 \$13246 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$42307 \$16 \$12032 \$16 \$153 \$13237 VNB sky130_fd_sc_hd__inv_1
X$42309 \$153 \$13291 \$12169 \$13207 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$42310 \$153 \$13290 \$12179 \$13237 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42312 \$153 \$13263 \$11881 \$13237 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42314 \$153 \$13016 \$12119 \$12907 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42315 \$153 \$13264 \$12182 \$13247 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42316 \$16 \$11945 \$16 \$153 \$13247 VNB sky130_fd_sc_hd__inv_1
X$42319 \$153 \$13292 \$11942 \$13247 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42320 \$153 \$13293 \$11881 \$13247 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42321 \$16 \$12384 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42322 \$153 \$11555 \$10376 \$11016 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42323 \$153 \$13208 \$13126 \$12120 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42324 \$153 \$13182 \$12179 \$13209 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42325 \$16 \$12120 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42328 \$153 \$13294 \$13156 \$12120 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42329 \$153 \$13210 \$12179 \$13248 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42330 \$153 \$13294 \$12182 \$13248 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42331 \$16 \$11798 \$16 \$153 \$13248 VNB sky130_fd_sc_hd__inv_1
X$42332 \$16 \$12120 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42333 \$153 \$13238 \$13265 \$12120 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42335 \$153 \$13238 \$12182 \$13249 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42336 \$16 \$11483 \$16 \$153 \$13249 VNB sky130_fd_sc_hd__inv_1
X$42337 \$16 \$12303 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42338 \$153 \$13211 \$13020 \$12303 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42339 \$153 \$12981 \$12371 \$12980 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42340 \$153 \$12827 \$12227 \$12980 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42341 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$42343 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$42344 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$42345 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$42346 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$42347 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$42350 \$153 \$13335 \$13213 \$12230 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42352 \$16 \$12158 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42353 \$16 \$11757 \$16 \$153 \$13336 VNB sky130_fd_sc_hd__inv_1
X$42354 \$153 \$13337 \$13213 \$12236 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42355 \$153 \$13338 \$13213 \$12003 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42356 \$16 \$12003 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42358 \$153 \$13266 \$12229 \$13336 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42360 \$16 \$11898 \$12779 \$13113 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$42361 \$153 \$13339 \$13130 \$12158 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42362 \$16 \$11898 \$16 \$153 \$13239 VNB sky130_fd_sc_hd__inv_1
X$42363 \$16 \$12158 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42364 \$153 \$13267 \$12229 \$13239 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42365 \$16 \$12093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42366 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$42369 \$153 \$13191 \$12412 \$12924 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42370 \$16 \$12236 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42371 \$153 \$13304 \$13250 \$12003 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42372 \$153 \$13304 \$11810 \$13369 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42373 \$16 \$12003 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42375 \$153 \$13340 \$13115 \$12230 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42378 \$153 \$13269 \$12057 \$13194 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42379 \$153 \$13131 \$11810 \$13194 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42380 \$16 \$12158 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42381 \$153 \$13326 \$11810 \$13215 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42382 \$153 \$13270 \$12057 \$13216 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42383 \$16 \$12093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42384 \$16 \$13215 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42385 \$153 \$13185 \$11810 \$13216 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42386 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$42389 \$153 \$13341 \$13272 \$12095 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42391 \$153 \$13342 \$13272 \$12093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42392 \$16 \$11485 \$16 \$153 \$13343 VNB sky130_fd_sc_hd__inv_1
X$42393 \$16 \$12093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42394 \$16 \$12003 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42395 \$153 \$13344 \$13305 \$12093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42397 \$16 \$11814 \$16 \$153 \$13215 VNB sky130_fd_sc_hd__inv_1
X$42398 \$16 \$11814 \$12897 \$13297 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$42399 \$153 \$13048 \$13305 \$12158 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42400 \$153 \$13298 \$11995 \$13273 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$42401 \$153 \$13306 \$11810 \$13108 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42402 \$153 \$13307 \$11810 \$13345 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42404 \$16 \$11995 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42406 \$16 \$12093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42407 \$153 \$13346 \$13298 \$12093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42409 \$16 \$11795 \$16 \$153 \$13345 VNB sky130_fd_sc_hd__inv_1
X$42411 \$153 \$13347 \$11949 \$13274 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$42412 \$153 \$13308 \$13118 \$12296 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42414 \$153 \$13308 \$12359 \$13105 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42415 \$16 \$12259 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42416 \$16 \$12296 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42417 \$16 \$11898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42418 \$153 \$13252 \$13118 \$12160 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42419 \$153 \$13348 \$13118 \$12101 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42420 \$153 \$13403 \$12476 \$13373 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42422 \$16 \$11757 \$16 \$153 \$13222 VNB sky130_fd_sc_hd__inv_1
X$42423 \$16 \$12101 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42424 \$153 \$13309 \$13220 \$12101 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42425 \$153 \$13309 \$12476 \$13222 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42426 \$153 \$13310 \$13275 \$12044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42427 \$153 \$13310 \$12068 \$13327 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42430 \$153 \$13388 \$13275 \$12083 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42432 \$153 \$13299 \$13276 \$12296 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42433 \$16 \$11721 \$16 \$153 \$13240 VNB sky130_fd_sc_hd__inv_1
X$42434 \$16 \$12296 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42435 \$16 \$11721 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42436 \$153 \$13311 \$13276 \$12083 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42438 \$153 \$13311 \$12174 \$13240 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42439 \$16 \$11485 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42440 \$16 \$11485 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42441 \$16 \$11485 \$16 \$153 \$13241 VNB sky130_fd_sc_hd__inv_1
X$42443 \$153 \$13278 \$13190 \$12044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42444 \$16 \$12044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42445 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$42446 \$16 \$11795 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42447 \$153 \$13328 \$12359 \$13241 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42449 \$16 \$11795 \$12785 \$13255 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$42451 \$153 \$13349 \$13224 \$12296 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42452 \$153 \$13350 \$13224 \$12044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42453 \$153 \$13256 \$13224 \$12101 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42455 \$16 \$11814 \$12785 \$13351 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$42456 \$16 \$12101 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42458 \$153 \$13280 \$12359 \$13051 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42459 \$16 \$12160 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42460 \$16 \$12101 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42461 \$153 \$13352 \$12999 \$12101 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42462 \$153 \$13312 \$12999 \$12241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42463 \$153 \$13312 \$12363 \$13077 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42464 \$16 \$12295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42466 \$153 \$13282 \$12155 \$13077 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42467 \$153 \$13329 \$12174 \$13243 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42468 \$16 \$12115 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42469 \$153 \$13313 \$13330 \$12115 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42470 \$153 \$13313 \$12234 \$13244 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42472 \$153 \$13331 \$12110 \$13244 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42475 \$16 \$12115 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42476 \$16 \$11374 \$16 \$153 \$13244 VNB sky130_fd_sc_hd__inv_1
X$42477 \$153 \$13314 \$13258 \$12115 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42478 \$153 \$13314 \$12234 \$13200 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42480 \$16 \$12326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42481 \$153 \$13353 \$13258 \$12326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42482 \$16 \$12115 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42483 \$16 \$11930 \$16 \$153 \$13200 VNB sky130_fd_sc_hd__inv_1
X$42486 \$153 \$13354 \$13315 \$12115 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42487 \$16 \$11930 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42489 \$16 \$12219 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42490 \$153 \$13301 \$13315 \$12219 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42491 \$16 \$11772 \$16 \$153 \$13245 VNB sky130_fd_sc_hd__inv_1
X$42492 \$153 \$13316 \$12198 \$13202 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$42494 \$153 \$13355 \$13316 \$12326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42495 \$16 \$12198 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42496 \$16 \$11772 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42497 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$42498 \$153 \$13317 \$12110 \$13302 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42499 \$153 \$13356 \$13285 \$12115 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42500 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$42501 \$16 \$12326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42503 \$153 \$13357 \$13285 \$12326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42504 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$42505 \$16 \$12164 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42506 \$153 \$13358 \$13054 \$12164 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42507 \$153 \$13204 \$12234 \$12648 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42509 \$153 \$13230 \$12309 \$12863 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42511 \$153 \$13359 \$13260 \$12115 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42512 \$153 \$13120 \$13260 \$12326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42514 \$16 \$12115 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42515 \$153 \$13318 \$13110 \$12115 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42516 \$16 \$11921 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42519 \$153 \$13318 \$12234 \$13205 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42521 \$16 \$12297 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42522 \$153 \$13288 \$13175 \$12297 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42523 \$16 \$12298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42525 \$16 \$11459 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42526 \$16 \$12164 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42527 \$153 \$13360 \$13175 \$12164 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42529 \$16 \$12326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42531 \$153 \$13319 \$13175 \$12326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42532 \$153 \$13319 \$12264 \$13149 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42534 \$153 \$13361 \$12918 \$11983 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42536 \$153 \$13332 \$11942 \$13362 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42537 \$16 \$11374 \$16 \$153 \$13362 VNB sky130_fd_sc_hd__inv_1
X$42540 \$153 \$13363 \$12918 \$12384 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42541 \$16 \$12384 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42542 \$16 \$12351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42544 \$16 \$12010 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42545 \$153 \$13364 \$13094 \$12010 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42546 \$153 \$13320 \$12179 \$13056 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42547 \$16 \$11930 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42549 \$16 \$12010 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42551 \$16 \$12384 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42554 \$153 \$13303 \$13152 \$12384 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42555 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$42557 \$16 \$11983 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42558 \$153 \$13206 \$13180 \$11983 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42559 \$153 \$13321 \$13180 \$12010 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42561 \$16 \$12010 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42562 \$16 \$12384 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42563 \$153 \$13333 \$12179 \$13181 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42564 \$153 \$13321 \$11942 \$13181 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42565 \$153 \$13290 \$13289 \$12384 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42566 \$153 \$13365 \$13289 \$12120 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42567 \$16 \$12120 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42569 \$153 \$13264 \$13291 \$12120 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42570 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$42571 \$16 \$11945 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42572 \$16 \$12384 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42573 \$153 \$13322 \$13291 \$12384 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42574 \$153 \$13322 \$12179 \$13247 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42575 \$16 \$11747 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42577 \$16 \$12010 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42578 \$16 \$12120 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42580 \$153 \$13323 \$13126 \$12010 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42581 \$153 \$13323 \$11942 \$13209 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42582 \$16 \$11459 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42583 \$16 \$11983 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42584 \$153 \$13324 \$13156 \$11983 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42586 \$153 \$13324 \$11881 \$13248 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42589 \$16 \$11776 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42590 \$16 \$11172 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42591 \$16 \$11798 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42592 \$16 \$12010 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42593 \$153 \$13334 \$12339 \$13248 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42594 \$153 \$13366 \$13265 \$12010 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42595 \$16 \$12782 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42596 \$16 \$11483 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42597 \$16 \$12384 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42598 \$153 \$13325 \$13265 \$12384 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42601 \$153 \$13325 \$12179 \$13249 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42602 \$153 \$12762 \$11881 \$12980 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42603 \$153 \$13025 \$12119 \$12980 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42604 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$42606 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$42607 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$42608 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$42609 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$42612 \$153 \$25 \$64 \$17 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42613 \$153 \$25 \$102 \$88 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42614 \$16 \$17 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42617 \$153 \$127 \$64 \$184 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42618 \$16 \$184 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42620 \$153 \$90 \$30 \$89 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42623 \$16 \$58 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42625 \$153 \$26 \$65 \$17 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42626 \$16 \$17 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42627 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$42629 \$153 \$26 \$102 \$89 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42631 \$153 \$91 \$59 \$94 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42632 \$153 \$92 \$377 \$94 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42634 \$153 \$93 \$102 \$94 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42635 \$16 \$17 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42637 \$153 \$128 \$66 \$17 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42640 \$153 \$95 \$30 \$96 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42641 \$16 \$17 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42642 \$153 \$129 \$67 \$58 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42644 \$16 \$58 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42646 \$153 \$97 \$102 \$270 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42647 \$153 \$130 \$68 \$184 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42649 \$153 \$131 \$68 \$17 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42650 \$153 \$130 \$59 \$98 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42651 \$16 \$17 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42655 \$16 \$58 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42656 \$153 \$99 \$59 \$100 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42657 \$153 \$27 \$190 \$17 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42659 \$153 \$27 \$102 \$100 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42660 \$16 \$17 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42661 \$153 \$28 \$69 \$17 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42664 \$153 \$28 \$102 \$101 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42665 \$16 \$17 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42667 \$153 \$132 \$70 \$17 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42669 \$16 \$17 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42670 \$153 \$29 \$70 \$58 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42671 \$153 \$29 \$30 \$172 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42674 \$153 \$103 \$59 \$172 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42676 \$16 \$58 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42677 \$153 \$31 \$71 \$58 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42679 \$16 \$17 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42681 \$153 \$31 \$30 \$173 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42682 \$153 \$32 \$72 \$187 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42684 \$16 \$187 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42686 \$153 \$32 \$54 \$174 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42687 \$153 \$133 \$72 \$73 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42689 \$16 \$73 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42690 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$42691 \$153 \$33 \$72 \$60 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42692 \$16 \$60 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42695 \$153 \$33 \$104 \$174 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42697 \$153 \$134 \$74 \$60 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42698 \$16 \$60 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42700 \$153 \$135 \$74 \$73 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42701 \$16 \$73 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42703 \$153 \$52 \$215 \$105 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42705 \$153 \$34 \$185 \$18 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42706 \$153 \$106 \$35 \$105 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42707 \$16 \$18 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42710 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$42711 \$153 \$136 \$24 \$18 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42713 \$16 \$18 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42714 \$16 \$18 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42715 \$153 \$137 \$24 \$60 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42716 \$16 \$60 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42717 \$16 \$73 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42718 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$42720 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$42721 \$153 \$138 \$53 \$73 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42722 \$16 \$60 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42723 \$16 \$73 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42724 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$42726 \$153 \$36 \$53 \$18 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42727 \$16 \$18 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42730 \$153 \$37 \$193 \$60 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42731 \$153 \$37 \$104 \$20 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42732 \$16 \$60 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42735 \$153 \$19 \$54 \$20 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42736 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$42737 \$153 \$139 \$194 \$73 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42739 \$16 \$60 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42740 \$153 \$38 \$75 \$60 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42743 \$153 \$38 \$104 \$329 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42744 \$16 \$73 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42745 \$153 \$39 \$75 \$73 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42748 \$153 \$39 \$215 \$329 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42750 \$16 \$79 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42753 \$153 \$140 \$76 \$79 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42756 \$153 \$109 \$44 \$352 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42757 \$16 \$79 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42758 \$153 \$141 \$61 \$79 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42761 \$153 \$110 \$44 \$111 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42763 \$16 \$82 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42764 \$153 \$55 \$112 \$113 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42765 \$153 \$55 \$77 \$79 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42769 \$153 \$114 \$559 \$113 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42772 \$153 \$41 \$559 \$115 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42775 \$153 \$56 \$112 \$177 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42777 \$16 \$591 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42779 \$16 \$80 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42780 \$16 \$79 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42781 \$153 \$56 \$267 \$79 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42783 \$16 \$116 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42786 \$16 \$145 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42787 \$153 \$118 \$21 \$117 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42789 \$153 \$43 \$81 \$82 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42790 \$153 \$43 \$44 \$117 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42791 \$16 \$80 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42794 \$153 \$119 \$266 \$117 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42795 \$16 \$82 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42796 \$153 \$146 \$62 \$82 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42799 \$153 \$146 \$44 \$120 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42800 \$16 \$145 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42803 \$153 \$45 \$21 \$120 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42806 \$153 \$46 \$23 \$121 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42807 \$16 \$178 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42810 \$153 \$47 \$83 \$63 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42811 \$153 \$47 \$57 \$121 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42814 \$153 \$22 \$84 \$310 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42815 \$16 \$310 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42817 \$153 \$123 \$398 \$122 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42819 \$153 \$48 \$85 \$310 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42820 \$153 \$48 \$223 \$122 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42824 \$153 \$125 \$23 \$124 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42826 \$16 \$399 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42827 \$16 \$258 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42828 \$16 \$258 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42829 \$16 \$63 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42830 \$153 \$49 \$227 \$63 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42831 \$16 \$149 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42833 \$153 \$49 \$57 \$124 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42836 \$16 \$151 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42837 \$16 \$63 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42838 \$16 \$149 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42839 \$16 \$63 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42842 \$16 \$178 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42844 \$16 \$80 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42845 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$42847 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$42848 \$16 \$63 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42849 \$153 \$201 \$50 \$63 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42850 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$42852 \$16 \$149 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42853 \$153 \$51 \$50 \$149 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42855 \$153 \$51 \$398 \$126 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42857 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$42859 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$42860 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$42861 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$42863 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$42865 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$42866 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$42867 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$42870 \$153 \$10861 \$10729 \$10368 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42871 \$153 \$10758 \$10729 \$10295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42872 \$16 \$10295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42873 \$16 \$10368 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42874 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$42875 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$42876 \$153 \$10662 \$10729 \$10200 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42878 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$42879 \$153 \$10903 \$10729 \$10367 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42880 \$153 \$10861 \$10303 \$10511 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42881 \$16 \$10367 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42882 \$16 \$10646 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42883 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$42884 \$16 \$10200 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42887 \$153 \$10759 \$10729 \$10476 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42888 \$153 \$10742 \$10729 \$10226 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42889 \$153 \$10904 \$10161 \$11055 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42890 \$153 \$10759 \$10705 \$10511 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42891 \$16 \$10764 \$16 \$153 \$10511 VNB sky130_fd_sc_hd__inv_1
X$42892 \$16 \$10764 \$10468 \$10842 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$42894 \$16 \$10226 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42895 \$16 \$10427 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42896 \$16 \$10888 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42897 \$153 \$10743 \$10594 \$10427 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42898 \$153 \$10862 \$10594 \$10476 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42899 \$16 \$10646 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42900 \$16 \$10476 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42901 \$16 \$10764 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42902 \$153 \$10905 \$10276 \$10884 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42903 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$42906 \$153 \$10843 \$10594 \$10367 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42907 \$153 \$10862 \$10705 \$10599 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42909 \$153 \$10843 \$10330 \$10599 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42910 \$16 \$10367 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42911 \$16 \$10744 \$16 \$153 \$10599 VNB sky130_fd_sc_hd__inv_1
X$42913 \$16 \$10427 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42914 \$16 \$10744 \$10468 \$10875 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$42915 \$153 \$10760 \$10532 \$10427 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42917 \$153 \$10594 \$10890 \$10875 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$42918 \$153 \$10760 \$10327 \$10745 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42919 \$153 \$10816 \$10532 \$10476 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42920 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$42921 \$16 \$10476 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42923 \$153 \$10816 \$10705 \$10745 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42924 \$153 \$10761 \$10276 \$10745 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42925 \$16 \$10427 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42927 \$153 \$10844 \$10652 \$10427 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42928 \$153 \$10906 \$10652 \$10226 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42929 \$153 \$10763 \$10652 \$10476 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42931 \$153 \$10844 \$10327 \$10746 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42932 \$153 \$10906 \$10161 \$10746 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42933 \$153 \$10763 \$10705 \$10746 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42935 \$153 \$10721 \$10652 \$10367 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42936 \$16 \$10476 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42937 \$16 \$10555 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42939 \$153 \$10765 \$10652 \$10368 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42940 \$16 \$10368 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42941 \$16 \$10825 \$10635 \$10876 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$42942 \$153 \$10652 \$11993 \$10876 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$42943 \$153 \$10765 \$10303 \$10746 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42944 \$16 \$10825 \$16 \$153 \$10746 VNB sky130_fd_sc_hd__inv_1
X$42946 \$153 \$10766 \$10524 \$10427 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42947 \$153 \$10863 \$10524 \$10476 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42948 \$153 \$10766 \$10327 \$10513 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42949 \$153 \$10863 \$10705 \$10513 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42951 \$16 \$10367 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42952 \$153 \$10707 \$10161 \$10513 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42954 \$153 \$10767 \$10524 \$10367 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42956 \$16 \$10747 \$16 \$153 \$10513 VNB sky130_fd_sc_hd__inv_1
X$42957 \$153 \$10524 \$10624 \$10748 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$42958 \$153 \$10767 \$10330 \$10513 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42959 \$16 \$10476 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42961 \$153 \$10768 \$10817 \$10226 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42962 \$16 \$10367 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42964 \$153 \$10864 \$10817 \$10367 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42965 \$153 \$10768 \$10161 \$10805 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42966 \$153 \$10864 \$10330 \$10805 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42967 \$16 \$10732 \$10635 \$10818 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$42968 \$153 \$10819 \$10817 \$10646 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42970 \$153 \$10456 \$10682 \$10818 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$42971 \$16 \$10732 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42972 \$153 \$10819 \$10318 \$10805 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42974 \$16 \$10200 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42976 \$153 \$10877 \$10907 \$10865 \$10885 \$10878 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$42978 \$153 \$153 \$10318 \$10602 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$42981 \$16 \$10886 \$16 \$153 \$10539 VNB sky130_fd_sc_hd__clkbuf_2
X$42982 \$16 \$10820 \$16 \$153 \$10348 VNB sky130_fd_sc_hd__clkbuf_2
X$42983 \$153 \$10887 \$10885 \$10877 \$10907 \$10878 \$16 \$16 VNB
+ sky130_fd_sc_hd__nor4b_2
X$42984 \$16 \$10295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42985 \$16 \$10634 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42986 \$153 \$10653 \$10634 \$10806 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$42987 \$16 \$10887 \$16 \$153 \$10453 VNB sky130_fd_sc_hd__clkbuf_2
X$42989 \$16 \$10888 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42990 \$153 \$10822 \$10888 \$10908 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$42992 \$16 \$10730 \$10525 \$10806 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$42993 \$16 \$10764 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42994 \$16 \$10730 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42995 \$16 \$10606 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42996 \$153 \$10910 \$10821 \$10526 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42997 \$153 \$10769 \$10821 \$10606 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$42998 \$16 \$10526 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$42999 \$16 \$10606 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43001 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$43002 \$153 \$10909 \$10538 \$10941 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43003 \$153 \$10771 \$10822 \$10338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43004 \$153 \$10709 \$10344 \$10477 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43006 \$16 \$10338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43007 \$153 \$10866 \$10822 \$10470 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43008 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$43011 \$153 \$10771 \$10309 \$10750 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43012 \$153 \$10889 \$10098 \$10941 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43013 \$153 \$10749 \$10822 \$10606 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43014 \$153 \$10866 \$10247 \$10750 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43015 \$16 \$10606 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43016 \$16 \$10470 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43019 \$153 \$10823 \$10822 \$10298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43020 \$153 \$10751 \$10822 \$10382 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43021 \$16 \$10382 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43022 \$153 \$10823 \$10401 \$10750 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43023 \$16 \$10890 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43024 \$153 \$10670 \$10890 \$10943 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$43025 \$16 \$10298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43027 \$153 \$10772 \$10670 \$10338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43028 \$153 \$10867 \$10670 \$10526 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43029 \$16 \$10338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43030 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$43031 \$153 \$10867 \$10516 \$10647 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43032 \$16 \$10744 \$16 \$153 \$10647 VNB sky130_fd_sc_hd__inv_1
X$43033 \$16 \$10526 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43036 \$16 \$10744 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43037 \$153 \$10824 \$10670 \$10298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43039 \$153 \$10911 \$10670 \$10605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43040 \$153 \$10772 \$10309 \$10647 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43041 \$16 \$10605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43042 \$16 \$10825 \$10655 \$10879 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$43043 \$153 \$10731 \$11993 \$10879 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$43046 \$153 \$10824 \$10401 \$10647 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43047 \$16 \$10825 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43049 \$153 \$10912 \$10731 \$10338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43050 \$153 \$10845 \$10731 \$10514 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43052 \$153 \$10685 \$10686 \$10515 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43054 \$153 \$10845 \$10538 \$10891 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43055 \$16 \$10514 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43056 \$16 \$10825 \$16 \$153 \$10891 VNB sky130_fd_sc_hd__inv_1
X$43057 \$153 \$10774 \$10731 \$10470 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43058 \$16 \$10338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43060 \$153 \$10868 \$10731 \$10526 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43062 \$153 \$10775 \$10731 \$10298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43063 \$16 \$10526 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43064 \$153 \$10868 \$10516 \$10891 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43065 \$153 \$10711 \$10098 \$10891 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43066 \$153 \$10775 \$10401 \$10891 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43067 \$16 \$10298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43069 \$16 \$10732 \$10655 \$10776 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$43070 \$16 \$10732 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43072 \$16 \$10747 \$10655 \$10869 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$43073 \$153 \$10041 \$8651 \$9845 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43074 \$16 \$10413 \$10655 \$10913 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$43075 \$16 \$10747 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43076 \$153 \$10826 \$10323 \$10605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43077 \$153 \$10915 \$10893 \$10526 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43079 \$153 \$10914 \$10247 \$10892 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43080 \$16 \$10605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43081 \$16 \$10747 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43082 \$153 \$10777 \$10344 \$10343 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43083 \$16 \$10526 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43085 \$153 \$10916 \$10893 \$10382 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43086 \$153 \$10826 \$10686 \$10343 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43087 \$16 \$10732 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43088 \$153 \$10687 \$10344 \$10608 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43090 \$16 \$10382 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43092 \$16 \$10606 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43093 \$16 \$10605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43095 \$16 \$10382 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43097 \$153 \$10807 \$10607 \$10526 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43098 \$153 \$10870 \$10607 \$10605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43099 \$16 \$10526 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43100 \$153 \$10870 \$10686 \$10608 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43103 \$153 \$10807 \$10516 \$10608 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43104 \$153 \$10945 \$10098 \$10894 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43106 \$16 \$10538 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43107 \$16 \$10527 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43108 \$153 \$153 \$10098 \$10753 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43109 \$16 \$10338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43111 \$16 \$7829 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43112 \$153 \$10895 \$10501 \$10609 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43113 \$16 \$16 \$153 VNB sky130_fd_sc_hd__conb_1
X$43115 \$153 \$153 \$10309 \$10753 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43118 \$153 \$10896 \$10309 \$10894 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43119 \$153 \$153 \$10247 \$10753 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43120 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$43121 \$16 \$10735 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43122 \$153 \$10827 \$10733 \$10735 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43123 \$16 \$9845 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43124 \$153 \$10827 \$10919 \$10609 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43126 \$16 \$7994 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43127 \$16 \$10809 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43128 \$153 \$10828 \$10919 \$11207 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43129 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$43130 \$16 \$11207 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43131 \$16 \$10611 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43132 \$153 \$10830 \$10733 \$10578 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43133 \$16 \$10300 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43134 \$153 \$10846 \$10733 \$10611 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43136 \$16 \$10578 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43137 \$16 \$10386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43139 \$153 \$10829 \$10833 \$11207 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43140 \$153 \$10733 \$12406 \$10917 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$43141 \$153 \$10808 \$10471 \$10609 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43142 \$153 \$10918 \$10734 \$10578 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43143 \$16 \$10831 \$16 \$153 \$10609 VNB sky130_fd_sc_hd__inv_1
X$43144 \$16 \$10578 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43147 \$153 \$10830 \$10370 \$10609 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43148 \$16 \$10833 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43149 \$16 \$10473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43150 \$16 \$10300 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43151 \$153 \$10612 \$10734 \$10473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43152 \$153 \$10778 \$10734 \$10300 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43153 \$16 \$12406 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43154 \$16 \$11207 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43156 \$153 \$10918 \$10370 \$10480 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43157 \$16 \$10831 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43159 \$16 \$10809 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43160 \$153 \$10596 \$10463 \$10809 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43161 \$153 \$10778 \$10417 \$10480 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43163 \$16 \$10809 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43164 \$16 \$10739 \$11127 \$10880 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$43165 \$16 \$10854 \$11127 \$10779 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$43166 \$153 \$10528 \$10897 \$10880 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$43168 \$153 \$10832 \$10833 \$10810 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43169 \$16 \$10735 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43170 \$153 \$10847 \$10528 \$10735 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43171 \$153 \$10756 \$10528 \$10809 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43172 \$16 \$10551 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43174 \$16 \$10611 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43175 \$153 \$10847 \$10919 \$10482 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43176 \$16 \$10739 \$16 \$153 \$10482 VNB sky130_fd_sc_hd__inv_1
X$43178 \$153 \$10848 \$10881 \$10611 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43179 \$16 \$10897 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43180 \$16 \$10739 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43181 \$16 \$10735 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43182 \$153 \$10920 \$10881 \$10735 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43183 \$16 \$10551 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43184 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$43186 \$16 \$10611 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43187 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$43188 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$43189 \$153 \$10781 \$10471 \$10373 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43190 \$16 \$10661 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43191 \$16 \$10300 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43192 \$153 \$10871 \$10882 \$10300 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43193 \$153 \$10689 \$10714 \$10373 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43194 \$16 \$12220 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43195 \$16 \$10736 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43196 \$153 \$10474 \$12220 \$10725 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$43198 \$153 \$10672 \$10833 \$10373 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43199 \$16 \$10735 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43200 \$16 \$10661 \$10737 \$10921 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$43201 \$153 \$10782 \$10404 \$10735 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43203 \$153 \$10922 \$10882 \$10473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43205 \$153 \$11042 \$10833 \$10811 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43206 \$153 \$10404 \$10615 \$10849 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$43207 \$16 \$10552 \$10737 \$10849 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$43208 \$153 \$10850 \$10834 \$10578 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43209 \$153 \$10715 \$10714 \$10757 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43211 \$153 \$10553 \$10833 \$10374 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43212 \$153 \$10851 \$10834 \$10611 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43213 \$153 \$10850 \$10370 \$10923 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43214 \$153 \$10851 \$10833 \$10923 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43215 \$153 \$10924 \$10834 \$10473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43218 \$153 \$10784 \$10475 \$10551 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43219 \$16 \$10551 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43220 \$16 \$10853 \$10737 \$10883 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$43221 \$153 \$10475 \$10852 \$10883 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$43222 \$153 \$10784 \$10471 \$10517 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43223 \$153 \$10783 \$10714 \$10517 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43226 \$153 \$10925 \$10658 \$10386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43227 \$153 \$10504 \$10472 \$10517 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43228 \$153 \$10442 \$10501 \$10517 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43229 \$153 \$10786 \$10370 \$10926 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43230 \$16 \$10852 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43231 \$16 \$10853 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43232 \$153 \$10925 \$10472 \$10926 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43235 \$153 \$10388 \$10860 \$10738 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$43236 \$16 \$10551 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43237 \$153 \$10927 \$10658 \$10300 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43238 \$153 \$10788 \$10658 \$10551 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43240 \$16 \$10409 \$16 \$153 \$10926 VNB sky130_fd_sc_hd__inv_1
X$43242 \$153 \$10787 \$10714 \$10926 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43243 \$153 \$10788 \$10471 \$10926 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43244 \$16 \$10898 \$16 \$153 \$10736 VNB sky130_fd_sc_hd__clkbuf_2
X$43245 \$16 \$10409 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43246 \$153 \$7091 \$8391 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$43247 \$16 \$10835 \$16 \$153 \$10661 VNB sky130_fd_sc_hd__clkbuf_2
X$43248 \$16 \$10478 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43249 \$16 \$10478 \$16 \$153 \$10648 VNB sky130_fd_sc_hd__clkbuf_2
X$43250 \$16 \$10836 \$16 \$153 \$10649 VNB sky130_fd_sc_hd__clkbuf_2
X$43253 \$16 \$10854 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43254 \$16 \$10854 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43255 \$16 \$10899 \$16 \$153 \$10597 VNB sky130_fd_sc_hd__clkbuf_2
X$43256 \$16 \$7091 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43257 \$153 \$10616 \$10780 \$10837 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$43258 \$16 \$10854 \$10838 \$10837 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$43259 \$16 \$10928 \$16 \$153 \$10529 VNB sky130_fd_sc_hd__clkbuf_2
X$43260 \$16 \$10900 \$16 \$153 \$10853 VNB sky130_fd_sc_hd__clkbuf_2
X$43261 \$16 \$10978 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43262 \$16 \$10929 \$16 \$153 \$10409 VNB sky130_fd_sc_hd__clkbuf_2
X$43263 \$16 \$10780 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43264 \$16 \$10854 \$16 \$153 \$10484 VNB sky130_fd_sc_hd__inv_1
X$43265 \$16 \$10564 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43267 \$153 \$10855 \$10839 \$10326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43268 \$153 \$10930 \$10839 \$10564 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43269 \$153 \$10855 \$10466 \$10812 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43271 \$153 \$10931 \$10839 \$10467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43272 \$16 \$10326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43275 \$153 \$10530 \$12406 \$10813 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$43276 \$16 \$10467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43277 \$16 \$12406 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43278 \$153 \$10932 \$10839 \$10446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43279 \$16 \$10831 \$10838 \$10813 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$43281 \$153 \$10856 \$10839 \$10393 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43282 \$16 \$10446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43285 \$16 \$10393 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43286 \$16 \$10617 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43287 \$153 \$10856 \$10694 \$10812 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43288 \$153 \$10857 \$10839 \$10346 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43289 \$153 \$10789 \$10376 \$10518 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43290 \$153 \$10857 \$10285 \$10812 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43291 \$16 \$10831 \$16 \$153 \$10518 VNB sky130_fd_sc_hd__inv_1
X$43294 \$16 \$10739 \$10838 \$10840 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$43296 \$153 \$10933 \$10740 \$10392 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43297 \$153 \$10444 \$10897 \$10840 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$43298 \$153 \$10674 \$10466 \$10518 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43299 \$16 \$9550 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43300 \$16 \$10392 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43301 \$16 \$10831 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43302 \$16 \$10393 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43304 \$153 \$10791 \$10740 \$10393 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43305 \$153 \$10872 \$10740 \$10446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43306 \$153 \$10791 \$10694 \$10814 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43307 \$153 \$10872 \$10376 \$10814 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43308 \$16 \$10739 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43309 \$16 \$10446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43312 \$16 \$10564 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43313 \$153 \$10792 \$10466 \$10814 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43314 \$153 \$10873 \$10901 \$10564 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43315 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$43316 \$16 \$12220 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43317 \$153 \$10394 \$12220 \$10793 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$43318 \$153 \$10873 \$10642 \$10902 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43319 \$16 \$10392 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43321 \$153 \$10874 \$10901 \$10392 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43322 \$153 \$10676 \$10815 \$10519 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43323 \$16 \$10736 \$16 \$153 \$10520 VNB sky130_fd_sc_hd__inv_1
X$43325 \$153 \$10395 \$12050 \$10677 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$43326 \$153 \$10874 \$10815 \$10902 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43327 \$16 \$10467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43329 \$16 \$10617 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43331 \$153 \$10934 \$10395 \$10467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43332 \$16 \$10649 \$16 \$153 \$10858 VNB sky130_fd_sc_hd__inv_1
X$43333 \$153 \$10859 \$10395 \$10617 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43334 \$16 \$10446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43335 \$153 \$10699 \$10587 \$10650 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43336 \$153 \$10325 \$10981 \$10698 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$43339 \$16 \$10392 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43340 \$16 \$10326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43341 \$153 \$10935 \$10995 \$10326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43342 \$16 \$10661 \$16 \$153 \$10650 VNB sky130_fd_sc_hd__inv_1
X$43343 \$153 \$10794 \$10325 \$10392 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43345 \$16 \$12245 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43346 \$153 \$10678 \$10815 \$10521 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43348 \$16 \$10346 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43350 \$16 \$10597 \$10644 \$10795 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$43351 \$153 \$10591 \$10587 \$10521 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43353 \$153 \$10700 \$10560 \$10521 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43354 \$153 \$10397 \$10960 \$10630 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$43355 \$153 \$10798 \$10796 \$10346 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43357 \$153 \$9781 \$8996 \$10222 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43358 \$16 \$10529 \$10644 \$10797 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$43359 \$16 \$10222 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43361 \$153 \$10936 \$10796 \$10393 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43362 \$153 \$10799 \$10592 \$10346 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43364 \$16 \$10564 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43367 \$153 \$10841 \$10796 \$10564 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43369 \$153 \$9783 \$9122 \$10510 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43370 \$153 \$9922 \$9059 \$10510 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43371 \$16 \$10510 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43373 \$153 \$9863 \$8923 \$10510 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43374 \$16 \$8102 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43375 \$153 \$8102 \$7463 \$7033 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43378 \$153 \$10937 \$10796 \$10617 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43380 \$153 \$10803 \$10592 \$10467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43381 \$16 \$7033 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43382 \$153 \$8103 \$7639 \$7033 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43384 \$16 \$7033 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43385 \$153 \$8254 \$7607 \$7033 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43387 \$16 \$8103 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43388 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$43389 \$16 \$8254 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43390 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$43391 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$43392 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$43393 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$43396 \$153 \$10255 \$10554 \$10295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43397 \$153 \$10531 \$10729 \$10427 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43398 \$16 \$10427 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43399 \$16 \$10295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43400 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$43401 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$43403 \$153 \$10030 \$10554 \$10200 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43405 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$43406 \$153 \$10703 \$10729 \$10646 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43407 \$153 \$10662 \$10088 \$10511 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43408 \$153 \$10703 \$10318 \$10511 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43409 \$16 \$10200 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43413 \$153 \$10758 \$10276 \$10511 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43414 \$153 \$10663 \$10554 \$10226 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43416 \$16 \$10476 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43417 \$153 \$10742 \$10161 \$10511 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43418 \$153 \$10554 \$10634 \$10651 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$43419 \$16 \$10730 \$10468 \$10651 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$43422 \$16 \$10764 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43423 \$153 \$10664 \$10594 \$10646 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43425 \$153 \$10593 \$10594 \$10295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43427 \$153 \$10743 \$10327 \$10599 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43428 \$16 \$10295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43429 \$16 \$10634 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43430 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$43432 \$153 \$10664 \$10318 \$10599 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43434 \$153 \$10704 \$10594 \$10226 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43435 \$153 \$10618 \$10088 \$10599 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43436 \$153 \$10704 \$10161 \$10599 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43437 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$43438 \$153 \$10665 \$10532 \$10367 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43439 \$16 \$10226 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43441 \$16 \$10744 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43442 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$43443 \$153 \$10533 \$10161 \$10745 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43444 \$16 \$10367 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43445 \$153 \$10619 \$10303 \$10745 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43446 \$153 \$10761 \$10532 \$10295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43447 \$16 \$10368 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43449 \$16 \$10523 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43451 \$153 \$10665 \$10330 \$10745 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43452 \$16 \$10295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43453 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$43454 \$16 \$10646 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43456 \$153 \$10679 \$10652 \$10200 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43457 \$153 \$10762 \$10652 \$10295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43458 \$16 \$10226 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43460 \$153 \$10679 \$10088 \$10746 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43461 \$16 \$10200 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43462 \$16 \$10295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43464 \$153 \$10720 \$10652 \$10646 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43465 \$153 \$10762 \$10276 \$10746 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43467 \$153 \$10720 \$10318 \$10746 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43468 \$16 \$10555 \$10635 \$10645 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$43470 \$16 \$10646 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43471 \$153 \$10259 \$10722 \$10645 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$43473 \$16 \$10476 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43474 \$153 \$10721 \$10330 \$10746 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43475 \$153 \$10620 \$10705 \$10212 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43476 \$153 \$10199 \$10706 \$10680 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$43477 \$16 \$10413 \$10635 \$10680 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$43480 \$153 \$10666 \$10524 \$10200 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43481 \$16 \$10413 \$16 \$153 \$10212 VNB sky130_fd_sc_hd__inv_1
X$43482 \$16 \$10427 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43483 \$16 \$10722 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43484 \$153 \$10707 \$10524 \$10226 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43485 \$153 \$10666 \$10088 \$10513 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43486 \$16 \$10226 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43487 \$16 \$10200 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43488 \$16 \$10825 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43489 \$16 \$10706 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43491 \$153 \$10600 \$10524 \$10646 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43492 \$16 \$10413 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43493 \$16 \$10747 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43494 \$16 \$10747 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43495 \$16 \$10747 \$10635 \$10748 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$43496 \$153 \$10252 \$10667 \$10681 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$43497 \$16 \$10621 \$10635 \$10681 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$43498 \$16 \$10646 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43499 \$16 \$10667 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43500 \$16 \$10427 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43501 \$16 \$10476 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43502 \$153 \$10636 \$10456 \$10427 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43504 \$153 \$10708 \$10456 \$10476 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43505 \$153 \$10636 \$10327 \$10334 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43506 \$153 \$10708 \$10705 \$10334 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43507 \$16 \$10732 \$16 \$153 \$10334 VNB sky130_fd_sc_hd__inv_1
X$43508 \$16 \$10646 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43511 \$153 \$10601 \$10456 \$10646 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43512 \$16 \$10682 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43513 \$16 \$10732 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43514 \$153 \$10683 \$10456 \$10368 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43515 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$43516 \$153 \$10683 \$10303 \$10334 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43517 \$16 \$10368 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43518 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$43519 \$153 \$153 \$10303 \$10602 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43521 \$153 \$153 \$10330 \$10602 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43522 \$16 \$16 \$153 VNB sky130_fd_sc_hd__conb_1
X$43525 \$153 \$153 \$10088 \$10602 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43526 \$153 \$153 \$10327 \$10602 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43528 \$16 \$10500 \$16 \$153 \$10602 VNB sky130_fd_sc_hd__clkbuf_2
X$43529 \$153 \$10709 \$10653 \$10606 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43530 \$16 \$10500 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43533 \$153 \$153 \$10161 \$10602 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43534 \$153 \$10669 \$10653 \$10526 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43535 \$153 \$10668 \$10653 \$10514 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43536 \$16 \$10514 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43537 \$16 \$10526 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43541 \$153 \$10770 \$10653 \$10605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43542 \$153 \$10669 \$10516 \$10477 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43543 \$153 \$10668 \$10538 \$10477 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43544 \$16 \$10605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43546 \$153 \$10654 \$10098 \$10477 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43547 \$16 \$10730 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43548 \$16 \$10730 \$16 \$153 \$10477 VNB sky130_fd_sc_hd__inv_1
X$43549 \$153 \$10654 \$10653 \$10382 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43551 \$153 \$10459 \$10653 \$10470 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43552 \$153 \$10622 \$10401 \$10477 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43553 \$153 \$10400 \$10522 \$10623 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$43554 \$16 \$10382 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43555 \$16 \$10470 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43557 \$16 \$10539 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43559 \$153 \$10749 \$10344 \$10750 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43560 \$16 \$10539 \$16 \$153 \$10337 VNB sky130_fd_sc_hd__inv_1
X$43562 \$153 \$10604 \$10400 \$10514 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43564 \$153 \$10751 \$10098 \$10750 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43565 \$153 \$10540 \$10686 \$10337 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43567 \$16 \$10453 \$10525 \$10541 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$43569 \$16 \$10514 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43570 \$16 \$10605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43572 \$16 \$10453 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43573 \$153 \$10637 \$10670 \$10514 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43574 \$153 \$10773 \$10670 \$10606 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43575 \$153 \$10637 \$10538 \$10647 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43576 \$16 \$10514 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43577 \$16 \$10606 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43578 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$43580 \$16 \$10453 \$16 \$153 \$10339 VNB sky130_fd_sc_hd__inv_1
X$43581 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$43582 \$16 \$10453 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43583 \$153 \$10710 \$10670 \$10470 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43585 \$153 \$10671 \$10670 \$10382 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43586 \$16 \$10298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43587 \$16 \$10470 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43588 \$16 \$10382 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43589 \$16 \$10722 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43591 \$16 \$10555 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43592 \$153 \$10381 \$10722 \$10684 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$43594 \$16 \$10555 \$10655 \$10684 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$43595 \$16 \$10605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43597 \$153 \$10685 \$10381 \$10605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43599 \$153 \$10723 \$10731 \$10605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43600 \$153 \$10710 \$10247 \$10647 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43602 \$153 \$10671 \$10098 \$10647 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43603 \$16 \$10621 \$10655 \$10656 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$43604 \$153 \$10752 \$10344 \$10891 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43605 \$153 \$10340 \$10667 \$10656 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$43606 \$16 \$10605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43607 \$16 \$10621 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43608 \$153 \$10711 \$10731 \$10382 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43609 \$16 \$10667 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43610 \$16 \$10621 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43612 \$16 \$10382 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43613 \$153 \$10545 \$10340 \$10606 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43614 \$153 \$10774 \$10247 \$10891 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43615 \$153 \$10546 \$10340 \$10514 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43616 \$153 \$10723 \$10686 \$10891 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43618 \$153 \$10607 \$10682 \$10776 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$43619 \$153 \$10323 \$10624 \$10869 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$43620 \$16 \$10682 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43621 \$153 \$10777 \$10323 \$10606 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43622 \$16 \$10514 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43623 \$16 \$10605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43624 \$16 \$9845 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43627 \$153 \$10625 \$10686 \$10249 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43628 \$16 \$10747 \$16 \$153 \$10343 VNB sky130_fd_sc_hd__inv_1
X$43629 \$16 \$10606 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43631 \$153 \$10712 \$10607 \$10298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43632 \$153 \$10687 \$10607 \$10606 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43633 \$16 \$10732 \$16 \$153 \$10608 VNB sky130_fd_sc_hd__inv_1
X$43634 \$16 \$10514 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43636 \$16 \$10298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43637 \$153 \$10712 \$10401 \$10608 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43638 \$16 \$10606 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43639 \$153 \$10638 \$10607 \$10382 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43640 \$153 \$9904 \$8277 \$9845 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43641 \$16 \$9845 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43642 \$16 \$10382 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43643 \$16 \$9845 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43645 \$16 \$7829 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43646 \$16 \$10470 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43647 \$16 \$10605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43648 \$16 \$10338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43650 \$16 \$9845 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43652 \$153 \$10638 \$10098 \$10608 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43653 \$16 \$10500 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43654 \$153 \$153 \$10344 \$10753 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43655 \$153 \$10558 \$10247 \$10608 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43656 \$153 \$153 \$10538 \$10753 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43657 \$16 \$10408 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43658 \$153 \$153 \$10401 \$10753 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43659 \$16 \$10500 \$16 \$153 \$10753 VNB sky130_fd_sc_hd__clkbuf_2
X$43661 \$16 \$10143 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43663 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43664 \$153 \$153 \$10516 \$10753 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43665 \$16 \$9339 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43667 \$153 \$10143 \$10809 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$43668 \$153 \$153 \$10686 \$10753 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43670 \$153 \$10610 \$10733 \$10809 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43671 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43673 \$153 \$10080 \$8340 \$10919 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43674 \$153 \$10755 \$10733 \$10300 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43676 \$153 \$9624 \$8917 \$8126 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43677 \$16 \$10919 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43679 \$16 \$8340 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43680 \$16 \$8126 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43681 \$153 \$10008 \$8340 \$10833 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43683 \$153 \$10724 \$10733 \$10386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43685 \$16 \$10386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43686 \$16 \$10611 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43687 \$153 \$10462 \$10734 \$10611 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43688 \$153 \$153 \$10833 \$10479 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43690 \$153 \$153 \$10919 \$10479 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43691 \$153 \$10755 \$10417 \$10609 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43692 \$153 \$153 \$10714 \$10479 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43693 \$153 \$10724 \$10472 \$10609 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43695 \$153 \$10613 \$10463 \$10551 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43696 \$16 \$10551 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43697 \$16 \$10735 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43699 \$153 \$10713 \$10463 \$10735 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43700 \$153 \$10614 \$10463 \$10611 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43701 \$153 \$10463 \$10780 \$10779 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$43702 \$16 \$10611 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43704 \$16 \$10854 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43707 \$153 \$10657 \$10833 \$10482 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43708 \$16 \$10854 \$16 \$153 \$10372 VNB sky130_fd_sc_hd__inv_1
X$43709 \$16 \$10780 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43710 \$16 \$10611 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43711 \$153 \$10657 \$10528 \$10611 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43712 \$153 \$10688 \$10528 \$10578 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43713 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$43714 \$16 \$10578 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43716 \$153 \$10550 \$10501 \$10482 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43717 \$153 \$10688 \$10370 \$10482 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43719 \$153 \$10756 \$10714 \$10482 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43720 \$16 \$10809 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43721 \$153 \$10689 \$10474 \$10809 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43723 \$153 \$10781 \$10474 \$10551 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43725 \$153 \$10672 \$10474 \$10611 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43726 \$16 \$10735 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43727 \$153 \$10673 \$10474 \$10735 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43729 \$16 \$10611 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43730 \$153 \$10673 \$10919 \$10373 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43731 \$16 \$10736 \$16 \$153 \$10373 VNB sky130_fd_sc_hd__inv_1
X$43733 \$153 \$10690 \$10404 \$10611 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43735 \$16 \$10809 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43736 \$16 \$10736 \$10737 \$10725 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$43737 \$153 \$10715 \$10404 \$10809 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43738 \$153 \$10502 \$10501 \$10373 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43739 \$16 \$10736 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43741 \$16 \$10809 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43744 \$153 \$10782 \$10919 \$10757 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43745 \$153 \$10580 \$10471 \$10757 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43746 \$153 \$10438 \$10370 \$10757 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43748 \$153 \$10691 \$10387 \$10809 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43749 \$16 \$10578 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43750 \$153 \$10691 \$10714 \$10374 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43751 \$153 \$10581 \$10471 \$10374 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43754 \$16 \$10597 \$10737 \$10726 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$43755 \$153 \$10387 \$12245 \$10726 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$43756 \$16 \$10611 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43758 \$16 \$10611 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43759 \$16 \$10809 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43760 \$153 \$10582 \$10919 \$10374 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43761 \$153 \$10783 \$10475 \$10809 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43762 \$16 \$10735 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43764 \$16 \$10578 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43766 \$153 \$10639 \$10475 \$10578 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43767 \$153 \$10785 \$10475 \$10611 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43768 \$153 \$10639 \$10370 \$10517 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43769 \$16 \$10853 \$16 \$153 \$10517 VNB sky130_fd_sc_hd__inv_1
X$43770 \$153 \$10692 \$10658 \$10611 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43773 \$153 \$10786 \$10658 \$10578 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43775 \$153 \$10584 \$10833 \$10375 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43776 \$16 \$10735 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43777 \$153 \$10693 \$10658 \$10735 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43778 \$16 \$10578 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43779 \$16 \$10611 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43783 \$16 \$10809 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43784 \$153 \$10585 \$10919 \$10375 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43785 \$16 \$10529 \$10737 \$10738 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$43787 \$153 \$10659 \$10388 \$10809 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43788 \$153 \$10787 \$10658 \$10809 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43790 \$153 \$10659 \$10714 \$10375 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43791 \$153 \$10693 \$10919 \$10926 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43793 \$16 \$10529 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43794 \$153 \$153 \$10815 \$10648 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43795 \$153 \$153 \$10466 \$10648 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43796 \$153 \$153 \$10587 \$10648 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43797 \$153 \$153 \$10560 \$10648 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43799 \$153 \$153 \$10642 \$10648 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43800 \$153 \$153 \$10694 \$10648 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43801 \$153 \$153 \$10285 \$10648 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43802 \$153 \$153 \$10376 \$10648 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43804 \$153 \$10716 \$10815 \$10484 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43805 \$153 \$10695 \$10616 \$10564 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43807 \$153 \$10716 \$10616 \$10392 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43808 \$16 \$10564 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43810 \$153 \$10588 \$10616 \$10467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43811 \$153 \$10695 \$10642 \$10484 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43812 \$16 \$10392 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43813 \$16 \$10467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43817 \$153 \$10717 \$10616 \$10393 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43818 \$153 \$10640 \$10616 \$10617 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43819 \$153 \$10717 \$10694 \$10484 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43820 \$153 \$10640 \$10560 \$10484 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43821 \$16 \$10393 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43822 \$16 \$10617 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43826 \$153 \$10789 \$10530 \$10446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43827 \$16 \$10617 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43828 \$153 \$10641 \$10530 \$10617 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43830 \$153 \$10790 \$10530 \$10392 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43831 \$153 \$10641 \$10560 \$10518 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43833 \$16 \$10346 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43834 \$153 \$10674 \$10530 \$10326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43835 \$153 \$10675 \$10530 \$10564 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43836 \$16 \$10326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43837 \$153 \$10675 \$10642 \$10518 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43838 \$16 \$10564 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43839 \$16 \$10326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43840 \$16 \$10739 \$16 \$153 \$10519 VNB sky130_fd_sc_hd__inv_1
X$43842 \$153 \$10676 \$10444 \$10392 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43843 \$153 \$10792 \$10740 \$10326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43845 \$16 \$10739 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43846 \$153 \$10626 \$10560 \$10519 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43848 \$16 \$10467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43849 \$16 \$10564 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43850 \$153 \$10718 \$10444 \$10467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43853 \$153 \$10643 \$10444 \$10564 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43854 \$153 \$10718 \$10587 \$10519 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43855 \$153 \$10643 \$10642 \$10519 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43856 \$16 \$10736 \$10644 \$10793 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$43858 \$16 \$10736 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43859 \$16 \$10736 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43861 \$16 \$10649 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43863 \$16 \$10392 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43864 \$16 \$10617 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43865 \$153 \$10719 \$10394 \$10392 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43866 \$153 \$10696 \$10394 \$10617 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43867 \$153 \$10696 \$10560 \$10520 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43868 \$16 \$10649 \$10644 \$10677 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$43869 \$16 \$12050 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43872 \$153 \$10627 \$10587 \$10520 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43874 \$16 \$10393 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43875 \$153 \$10697 \$10395 \$10393 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43876 \$153 \$10419 \$10466 \$10520 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43877 \$153 \$10719 \$10815 \$10520 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43878 \$16 \$10661 \$10644 \$10698 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$43880 \$16 \$10467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43881 \$16 \$10564 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43882 \$153 \$10629 \$10560 \$10650 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43884 \$153 \$10727 \$10642 \$10650 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43885 \$153 \$10699 \$10325 \$10467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43886 \$153 \$10727 \$10325 \$10564 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43887 \$16 \$10392 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43888 \$16 \$10617 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43889 \$153 \$10396 \$12245 \$10795 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$43891 \$153 \$9990 \$8923 \$10222 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43892 \$153 \$10678 \$10396 \$10392 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43893 \$16 \$10222 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43895 \$153 \$10592 \$10860 \$10797 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$43896 \$16 \$10597 \$16 \$153 \$10521 VNB sky130_fd_sc_hd__inv_1
X$43899 \$153 \$10700 \$10396 \$10617 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43900 \$16 \$8429 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43901 \$153 \$8775 \$7639 \$8429 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43902 \$153 \$10800 \$10592 \$10393 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43903 \$16 \$10564 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43904 \$153 \$9921 \$8996 \$10510 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43905 \$16 \$10529 \$16 \$153 \$10741 VNB sky130_fd_sc_hd__inv_1
X$43908 \$153 \$10701 \$10397 \$10564 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43909 \$16 \$10510 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43910 \$16 \$10409 \$16 \$153 \$10801 VNB sky130_fd_sc_hd__inv_1
X$43911 \$153 \$10802 \$10592 \$10326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43912 \$153 \$9647 \$9256 \$9646 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43914 \$16 \$10467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43915 \$16 \$10326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43916 \$16 \$10617 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43919 \$16 \$7033 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43920 \$16 \$10392 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43921 \$153 \$10702 \$10592 \$10392 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43922 \$153 \$10804 \$10592 \$10617 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43923 \$153 \$9830 \$9059 \$9646 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43924 \$16 \$10409 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43926 \$16 \$7033 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43927 \$153 \$10728 \$7376 \$7033 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43929 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$43930 \$16 \$10728 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43931 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$43932 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$43933 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$43934 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$43935 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$43936 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$43938 \$153 \$6538 \$6403 \$5403 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43940 \$153 \$6477 \$6403 \$5245 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43941 \$16 \$5403 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43942 \$16 \$5245 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43943 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$43944 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$43946 \$153 \$6539 \$6403 \$5736 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43947 \$153 \$6430 \$4706 \$6452 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43948 \$153 \$6430 \$6403 \$5274 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43949 \$16 \$5736 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43951 \$153 \$6352 \$5463 \$6174 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43954 \$153 \$6526 \$5177 \$6452 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43955 \$16 \$4902 \$16 \$153 \$6452 VNB sky130_fd_sc_hd__inv_1
X$43956 \$153 \$6478 \$6397 \$5736 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43957 \$153 \$6478 \$5055 \$6257 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43958 \$153 \$6517 \$5177 \$6257 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43959 \$16 \$5489 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43960 \$16 \$5274 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43961 \$153 \$6404 \$6397 \$5245 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43964 \$16 \$5736 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43965 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$43966 \$16 \$4893 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43967 \$153 \$6527 \$5174 \$6257 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43968 \$153 \$6258 \$6397 \$5403 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43969 \$16 \$5245 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43970 \$16 \$5314 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43971 \$16 \$4893 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43972 \$16 \$5403 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43973 \$153 \$6497 \$6251 \$5736 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43976 \$153 \$6405 \$6251 \$5404 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43977 \$153 \$6498 \$6406 \$5736 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43978 \$16 \$5404 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43979 \$16 \$5403 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43981 \$16 \$5736 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43982 \$153 \$6319 \$6406 \$5403 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43984 \$153 \$6497 \$5055 \$6260 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43986 \$153 \$6407 \$4706 \$6315 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43987 \$16 \$5404 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43989 \$153 \$6458 \$6406 \$5245 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$43990 \$16 \$5274 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43991 \$16 \$5403 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43993 \$16 \$4896 \$16 \$153 \$6315 VNB sky130_fd_sc_hd__inv_1
X$43995 \$153 \$6458 \$5107 \$6315 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$43996 \$16 \$5245 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43997 \$16 \$4896 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$43998 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$43999 \$153 \$6499 \$6398 \$5404 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44000 \$153 \$6479 \$5463 \$6315 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44001 \$153 \$6408 \$5107 \$6409 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44002 \$16 \$5404 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44003 \$16 \$5736 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44006 \$153 \$6431 \$6398 \$5403 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44007 \$16 \$4621 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44008 \$153 \$6500 \$6398 \$5518 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44009 \$153 \$6431 \$5405 \$6409 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44010 \$153 \$6500 \$5463 \$6409 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44011 \$16 \$5274 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44013 \$16 \$5403 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44015 \$153 \$6378 \$6280 \$5736 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44016 \$16 \$4973 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44018 \$153 \$6518 \$5463 \$6412 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44019 \$153 \$6410 \$5405 \$6412 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44020 \$16 \$5736 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44022 \$153 \$6411 \$6280 \$5274 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44023 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$44025 \$153 \$6460 \$6280 \$5245 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44026 \$153 \$6459 \$5177 \$6412 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44027 \$153 \$6460 \$5107 \$6412 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44028 \$16 \$5274 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44029 \$16 \$5245 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44030 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$44031 \$153 \$6501 \$6341 \$5404 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44034 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$44035 \$153 \$6480 \$6341 \$5403 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44036 \$153 \$6501 \$5177 \$6316 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44037 \$16 \$5403 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44038 \$16 \$5404 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44040 \$16 \$5245 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44041 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$44042 \$153 \$6481 \$6341 \$5245 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44045 \$16 \$3335 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44046 \$153 \$6481 \$5107 \$6316 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44047 \$153 \$6482 \$6341 \$5736 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44048 \$153 \$3335 \$5245 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$44050 \$153 \$6432 \$5405 \$6044 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44051 \$153 \$3276 \$5404 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$44052 \$16 \$3276 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44053 \$16 \$5403 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44054 \$16 \$5736 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44055 \$16 \$4822 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44056 \$16 \$5274 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44057 \$153 \$6433 \$6399 \$5274 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44058 \$16 \$5404 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44061 \$16 \$6695 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44063 \$16 \$5489 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44064 \$153 \$6519 \$5373 \$6177 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44065 \$153 \$6342 \$6399 \$5245 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44066 \$16 \$2414 \$16 \$153 \$6540 VNB sky130_fd_sc_hd__clkbuf_2
X$44067 \$16 \$2414 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44068 \$16 \$3244 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44069 \$16 \$5245 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44070 \$153 \$3244 \$5736 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$44071 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$44073 \$16 \$4822 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44074 \$16 \$4822 \$16 \$153 \$6177 VNB sky130_fd_sc_hd__inv_1
X$44075 \$153 \$6285 \$5055 \$6045 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44076 \$16 \$5736 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44077 \$153 \$6528 \$5174 \$6177 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44078 \$153 \$6461 \$5209 \$6453 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44079 \$16 \$4902 \$5900 \$6434 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$44080 \$153 \$6436 \$6435 \$5271 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44082 \$153 \$6461 \$6435 \$5338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44083 \$153 \$6436 \$5069 \$6453 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44084 \$16 \$5338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44085 \$16 \$5900 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44086 \$16 \$4902 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44087 \$16 \$5271 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44089 \$16 \$5226 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44090 \$153 \$6541 \$6435 \$5469 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44093 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$44094 \$153 \$6462 \$6353 \$5467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44095 \$153 \$6380 \$5096 \$6414 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44096 \$16 \$5467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44097 \$16 \$5469 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44099 \$153 \$6437 \$5287 \$6414 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44100 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$44102 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$44103 \$153 \$6438 \$6353 \$5232 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44105 \$153 \$6286 \$5209 \$6414 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44106 \$153 \$6415 \$5069 \$6414 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44107 \$153 \$6438 \$5205 \$6414 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44108 \$16 \$5478 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44110 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$44111 \$16 \$5232 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44112 \$153 \$6502 \$6287 \$5469 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44113 \$153 \$6439 \$6287 \$5467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44114 \$153 \$6439 \$5406 \$6262 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44115 \$153 \$6502 \$5287 \$6262 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44116 \$16 \$5469 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44119 \$153 \$6355 \$5519 \$6262 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44120 \$16 \$5467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44121 \$16 \$5566 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44122 \$16 \$4939 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44123 \$153 \$6463 \$6326 \$5467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44124 \$16 \$6695 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44126 \$153 \$6503 \$6326 \$5324 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44127 \$16 \$5467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44129 \$16 \$4893 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44131 \$153 \$6503 \$5096 \$6264 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44132 \$153 \$6356 \$5069 \$6264 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44133 \$16 \$5324 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44134 \$153 \$6464 \$5287 \$6264 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44136 \$153 \$6542 \$6440 \$5324 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44137 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$44138 \$153 \$6441 \$6440 \$5338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44141 \$153 \$6543 \$6440 \$5467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44142 \$153 \$6441 \$5209 \$6357 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44143 \$153 \$6529 \$5287 \$6357 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44144 \$16 \$5338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44145 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$44147 \$16 \$5467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44149 \$153 \$6504 \$6344 \$5469 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44150 \$153 \$6442 \$6344 \$5467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44151 \$153 \$6442 \$5406 \$6358 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44152 \$153 \$6504 \$5287 \$6358 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44153 \$16 \$5469 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44154 \$16 \$5467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44156 \$16 \$4947 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44159 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$44160 \$153 \$6530 \$5096 \$6358 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44161 \$153 \$6483 \$6001 \$5566 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44162 \$153 \$6505 \$6001 \$5469 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44163 \$16 \$5566 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44164 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$44166 \$153 \$6505 \$5287 \$6122 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44167 \$153 \$6454 \$6001 \$5324 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44168 \$16 \$5469 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44170 \$153 \$6531 \$5390 \$6122 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44171 \$153 \$6454 \$5096 \$6122 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44172 \$16 \$5478 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44173 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$44174 \$16 \$5324 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44175 \$153 \$6484 \$6034 \$5469 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44177 \$153 \$6506 \$6034 \$5324 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44178 \$153 \$6384 \$5406 \$6122 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44179 \$153 \$6506 \$5096 \$6291 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44180 \$16 \$5324 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44181 \$153 \$6484 \$5287 \$6291 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44182 \$16 \$5469 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44184 \$153 \$6345 \$6361 \$5467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44186 \$16 \$4822 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44187 \$153 \$6520 \$5390 \$6416 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44188 \$16 \$4822 \$16 \$153 \$6416 VNB sky130_fd_sc_hd__inv_1
X$44189 \$153 \$6465 \$6361 \$5271 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44190 \$153 \$6521 \$5287 \$6416 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44192 \$153 \$6521 \$6361 \$5469 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44193 \$153 \$6465 \$5069 \$6416 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44194 \$153 \$6417 \$5209 \$6416 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44195 \$153 \$3373 \$5324 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$44196 \$16 \$5271 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44199 \$153 \$3720 \$5338 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$44200 \$153 \$1775 \$5796 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$44201 \$153 \$6443 \$6265 \$5819 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44203 \$153 \$6507 \$6265 \$5796 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44204 \$153 \$6466 \$6265 \$5605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44205 \$153 \$6507 \$5775 \$6418 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44206 \$16 \$5605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44207 \$16 \$5796 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44208 \$16 \$5702 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44211 \$153 \$6466 \$5625 \$6418 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44212 \$153 \$6508 \$6265 \$5528 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44213 \$153 \$6467 \$5470 \$6418 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44214 \$153 \$6508 \$5500 \$6418 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44215 \$16 \$5351 \$6252 \$6485 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$44217 \$16 \$5605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44218 \$16 \$5528 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44219 \$16 \$5528 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44222 \$153 \$6444 \$6332 \$5528 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44223 \$153 \$6509 \$6332 \$5605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44224 \$153 \$6444 \$5500 \$6267 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44225 \$153 \$6509 \$5625 \$6267 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44227 \$16 \$5796 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44228 \$153 \$6544 \$6332 \$5702 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44230 \$153 \$6522 \$6332 \$5796 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44231 \$153 \$6522 \$5775 \$6267 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44232 \$16 \$4834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44233 \$16 \$4780 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44235 \$16 \$5528 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44237 \$16 \$5714 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44238 \$153 \$6445 \$6333 \$5528 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44240 \$16 \$5702 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44242 \$153 \$6545 \$6333 \$5702 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44243 \$153 \$6445 \$5500 \$6234 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44244 \$16 \$4949 \$6252 \$6510 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$44246 \$16 \$5605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44248 \$16 \$4949 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44249 \$153 \$6546 \$6333 \$5605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44251 \$16 \$5796 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44253 \$153 \$6419 \$6333 \$5796 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44254 \$16 \$4949 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44256 \$153 \$6511 \$5498 \$6523 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$44258 \$16 \$5498 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44259 \$16 \$5528 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44260 \$153 \$6446 \$6253 \$5528 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44262 \$16 \$5017 \$6252 \$6523 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$44263 \$153 \$6512 \$6511 \$5714 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44265 \$153 \$6446 \$5500 \$6421 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44266 \$16 \$5796 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44267 \$16 \$5017 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44268 \$153 \$6420 \$6253 \$5796 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44270 \$16 \$5819 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44272 \$153 \$6524 \$6253 \$5819 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44273 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$44274 \$153 \$6524 \$6200 \$6421 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44275 \$16 \$5353 \$6269 \$6468 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$44276 \$16 \$6269 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44277 \$153 \$6563 \$5473 \$6468 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$44278 \$16 \$5353 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44279 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$44281 \$153 \$6532 \$6200 \$6533 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44282 \$16 \$5473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44284 \$16 \$5605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44285 \$16 \$5353 \$16 \$153 \$6533 VNB sky130_fd_sc_hd__inv_1
X$44286 \$153 \$6486 \$6238 \$5605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44287 \$153 \$6422 \$6238 \$5796 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44289 \$16 \$5702 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44290 \$153 \$6547 \$6238 \$5702 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44292 \$16 \$5528 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44293 \$153 \$6525 \$6238 \$5528 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44295 \$153 \$6525 \$5500 \$6176 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44296 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$44297 \$16 \$5834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44298 \$16 \$5714 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44299 \$16 \$5528 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44301 \$153 \$6487 \$6400 \$5528 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44302 \$153 \$6548 \$6400 \$5714 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44303 \$153 \$6423 \$5881 \$6455 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44304 \$153 \$6487 \$5500 \$6455 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44305 \$16 \$5819 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44306 \$153 \$6534 \$5625 \$6455 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44309 \$16 \$5702 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44310 \$16 \$6269 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44311 \$153 \$6424 \$6200 \$6455 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44312 \$153 \$6548 \$5755 \$6455 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44313 \$153 \$6470 \$4831 \$6469 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$44314 \$16 \$5834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44315 \$16 \$5819 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44316 \$153 \$6489 \$5755 \$6535 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44317 \$153 \$6488 \$6470 \$5819 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44319 \$153 \$6549 \$6470 \$5834 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44320 \$16 \$5702 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44321 \$16 \$6269 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44322 \$153 \$6425 \$6470 \$5702 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44323 \$153 \$6366 \$5470 \$6318 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44325 \$16 \$4830 \$6269 \$6469 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$44326 \$153 \$6549 \$5881 \$6535 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44328 \$153 \$6489 \$6470 \$5714 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44329 \$16 \$5714 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44330 \$16 \$4831 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44331 \$16 \$1673 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44332 \$153 \$6536 \$5938 \$6273 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44333 \$16 \$5767 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44334 \$153 \$6471 \$5627 \$6273 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44336 \$16 \$4834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44338 \$153 \$6471 \$6349 \$5887 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44339 \$153 \$6490 \$6349 \$5767 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44341 \$16 \$5887 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44342 \$153 \$6490 \$5575 \$6273 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44343 \$16 \$4830 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44344 \$16 \$4830 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44347 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$44348 \$16 \$1544 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44350 \$16 \$5351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44351 \$153 \$6491 \$6349 \$5609 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44352 \$153 \$6472 \$6349 \$5963 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44353 \$153 \$6472 \$5806 \$6273 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44354 \$16 \$5963 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44355 \$16 \$5609 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44356 \$16 \$5786 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44358 \$16 \$5767 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44359 \$153 \$6550 \$6244 \$5786 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44361 \$153 \$6473 \$5074 \$6367 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44362 \$153 \$6447 \$5575 \$6367 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44363 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$44364 \$16 \$5636 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44366 \$153 \$6513 \$6244 \$5636 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44367 \$16 \$5259 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44368 \$16 \$5887 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44370 \$153 \$6448 \$6244 \$5887 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44371 \$153 \$6513 \$5509 \$6367 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44372 \$153 \$6448 \$5627 \$6367 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44373 \$153 \$5939 \$5627 \$5475 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44374 \$16 \$5963 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44375 \$16 \$5636 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44377 \$16 \$5718 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44378 \$153 \$6514 \$6206 \$5636 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44379 \$153 \$6090 \$5635 \$5475 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44380 \$153 \$6474 \$6206 \$5609 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44381 \$153 \$6514 \$5509 \$6047 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44382 \$16 \$5609 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44384 \$16 \$5767 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44385 \$16 \$5786 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44386 \$153 \$6515 \$6401 \$5767 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44387 \$153 \$6449 \$6401 \$5786 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44388 \$153 \$6515 \$5575 \$6456 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44389 \$153 \$6449 \$5635 \$6456 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44391 \$16 \$4949 \$16 \$153 \$6456 VNB sky130_fd_sc_hd__inv_1
X$44393 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$44394 \$16 \$4949 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44395 \$16 \$5887 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44396 \$16 \$5579 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44397 \$153 \$6426 \$6401 \$5887 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44398 \$153 \$6516 \$6401 \$5579 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44399 \$16 \$5400 \$6255 \$6492 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$44400 \$153 \$6516 \$5484 \$6456 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44404 \$16 \$4562 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44405 \$16 \$4609 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44406 \$16 \$5400 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44407 \$16 \$5579 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44408 \$16 \$5609 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44409 \$153 \$6551 \$6308 \$5609 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44410 \$153 \$6450 \$6308 \$5579 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44411 \$153 \$6450 \$5484 \$6311 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44412 \$16 \$5400 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44414 \$16 \$4562 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44416 \$16 \$5887 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44417 \$16 \$5767 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44418 \$16 \$5718 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44419 \$153 \$6475 \$6308 \$5767 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44420 \$153 \$6312 \$6308 \$5718 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44421 \$16 \$4837 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44423 \$153 \$6351 \$5473 \$6493 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$44424 \$16 \$5353 \$6255 \$6493 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$44426 \$153 \$6475 \$5575 \$6311 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44427 \$153 \$6552 \$6351 \$5609 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44428 \$16 \$5636 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44429 \$153 \$6494 \$6351 \$5636 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44430 \$16 \$5609 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44431 \$16 \$4963 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44432 \$16 \$5353 \$16 \$153 \$6924 VNB sky130_fd_sc_hd__inv_1
X$44434 \$16 \$4831 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44436 \$153 \$6495 \$6351 \$5963 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44437 \$16 \$5887 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44438 \$153 \$6553 \$6351 \$5887 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44439 \$153 \$6476 \$5938 \$6457 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44441 \$16 \$5354 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44442 \$153 \$6537 \$5806 \$6457 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44444 \$16 \$4830 \$6255 \$6600 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$44445 \$153 \$6554 \$6562 \$5767 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44446 \$16 \$5767 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44448 \$153 \$6428 \$6256 \$5963 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44449 \$16 \$4830 \$16 \$153 \$6457 VNB sky130_fd_sc_hd__inv_1
X$44450 \$16 \$4830 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44451 \$153 \$6371 \$5484 \$6274 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44452 \$16 \$4830 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44455 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$44456 \$16 \$5887 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44457 \$16 \$5636 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44458 \$153 \$6496 \$6256 \$5887 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44459 \$153 \$6555 \$6562 \$5636 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44460 \$153 \$6429 \$5509 \$6274 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44461 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$44464 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$44465 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$44466 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$44467 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$44468 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$44469 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$44470 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$44471 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$44473 \$153 \$5807 \$5710 \$5181 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44474 \$153 \$5728 \$5710 \$5245 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44475 \$16 \$5181 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44476 \$16 \$5245 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44477 \$16 \$5403 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44478 \$153 \$5728 \$5107 \$5762 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44480 \$153 \$5807 \$5174 \$5762 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44481 \$153 \$5693 \$5405 \$5762 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44482 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$44483 \$153 \$5836 \$5710 \$5489 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44484 \$153 \$5768 \$5055 \$5762 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44485 \$16 \$5518 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44488 \$16 \$5489 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44489 \$16 \$4320 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44490 \$16 \$5376 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44491 \$153 \$5729 \$4706 \$5762 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44492 \$16 \$4320 \$16 \$153 \$5837 VNB sky130_fd_sc_hd__inv_1
X$44493 \$153 \$5769 \$5710 \$5404 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44494 \$16 \$4162 \$5176 \$5730 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$44495 \$16 \$5176 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44497 \$153 \$5769 \$5177 \$5762 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44498 \$16 \$5404 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44499 \$16 \$5518 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44501 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$44502 \$16 \$4162 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44503 \$16 \$3638 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44505 \$153 \$5808 \$5628 \$5489 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44506 \$153 \$5790 \$5628 \$5518 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44508 \$153 \$5808 \$5373 \$5618 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44509 \$16 \$5518 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44512 \$153 \$5639 \$5628 \$5403 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44514 \$153 \$5838 \$5628 \$5245 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44515 \$16 \$5403 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44517 \$16 \$4179 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44518 \$153 \$5628 \$4179 \$5731 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$44519 \$16 \$5245 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44521 \$16 \$4178 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44523 \$16 \$4178 \$5712 \$5871 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$44525 \$16 \$4269 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44526 \$16 \$4178 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44527 \$153 \$5791 \$5641 \$5404 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44528 \$153 \$5770 \$5641 \$5403 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44529 \$153 \$5791 \$5177 \$5619 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44530 \$16 \$5404 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44533 \$153 \$5732 \$5641 \$5518 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44534 \$16 \$5403 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44535 \$16 \$4479 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44536 \$153 \$5763 \$5641 \$5736 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44537 \$16 \$5518 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44538 \$16 \$3879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44539 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$44540 \$153 \$5733 \$5174 \$5619 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44541 \$16 \$5736 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44544 \$16 \$5388 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44545 \$16 \$5181 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44546 \$153 \$5643 \$4706 \$5619 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44547 \$16 \$5720 \$16 \$153 \$6051 VNB sky130_fd_sc_hd__clkbuf_2
X$44548 \$153 \$5809 \$5711 \$5181 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44549 \$153 \$5770 \$5405 \$5619 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44551 \$16 \$5245 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44552 \$153 \$5809 \$5174 \$5721 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44555 \$153 \$5920 \$5055 \$5721 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44556 \$16 \$4106 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44557 \$153 \$5810 \$5711 \$5489 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44558 \$153 \$5763 \$5055 \$5619 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44559 \$16 \$5518 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44560 \$16 \$5720 \$16 \$153 \$5712 VNB sky130_fd_sc_hd__clkbuf_2
X$44561 \$16 \$4600 \$5712 \$5839 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$44562 \$153 \$5734 \$5405 \$5721 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44564 \$153 \$5810 \$5373 \$5721 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44565 \$16 \$4146 \$5712 \$5873 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$44566 \$16 \$5720 \$16 \$153 \$5630 VNB sky130_fd_sc_hd__clkbuf_2
X$44567 \$16 \$5489 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44569 \$153 \$5811 \$5645 \$5403 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44570 \$16 \$3198 \$16 \$153 \$5720 VNB sky130_fd_sc_hd__clkbuf_2
X$44572 \$153 \$5771 \$5055 \$5621 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44575 \$16 \$5403 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44576 \$153 \$5812 \$5645 \$5404 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44577 \$16 \$4146 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44578 \$153 \$5586 \$5373 \$5621 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44579 \$153 \$5811 \$5405 \$5621 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44580 \$153 \$5812 \$5177 \$5621 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44582 \$153 \$5647 \$5461 \$5403 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44583 \$16 \$5404 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44585 \$153 \$5813 \$5461 \$5736 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44587 \$16 \$4494 \$5630 \$5792 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$44588 \$153 \$5735 \$5174 \$5517 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44589 \$153 \$5813 \$5055 \$5517 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44590 \$153 \$5949 \$5107 \$5621 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44591 \$16 \$5736 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44593 \$153 \$5793 \$5461 \$5404 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44595 \$16 \$5274 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44596 \$153 \$5793 \$5177 \$5517 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44597 \$16 \$5404 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44600 \$153 \$5737 \$5466 \$5274 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44601 \$153 \$5950 \$4706 \$5722 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44603 \$153 \$5723 \$5832 \$5245 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44605 \$153 \$5738 \$5373 \$5464 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44606 \$153 \$5737 \$4706 \$5464 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44607 \$153 \$5840 \$5832 \$5403 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44608 \$16 \$3886 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44610 \$16 \$4494 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44611 \$153 \$5665 \$5405 \$5464 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44613 \$153 \$5589 \$5463 \$5464 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44614 \$16 \$4494 \$16 \$153 \$5722 VNB sky130_fd_sc_hd__inv_1
X$44615 \$153 \$5833 \$5376 \$5841 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$44616 \$16 \$5376 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44618 \$153 \$5764 \$5406 \$5564 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44619 \$153 \$5739 \$5548 \$5271 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44621 \$153 \$5842 \$5833 \$5338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44622 \$153 \$5739 \$5069 \$5622 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44623 \$153 \$5740 \$5209 \$5622 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44624 \$16 \$5271 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44625 \$16 \$5338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44628 \$153 \$5649 \$5096 \$5564 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44630 \$153 \$5724 \$5548 \$5232 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44631 \$153 \$5843 \$5833 \$5478 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44632 \$16 \$5232 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44633 \$153 \$5826 \$5520 \$5271 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44634 \$16 \$5478 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44635 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$44638 \$153 \$5826 \$5069 \$5564 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44639 \$153 \$5764 \$5520 \$5467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44640 \$153 \$5741 \$5390 \$5564 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44641 \$153 \$5844 \$5096 \$5845 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44642 \$16 \$5271 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44643 \$16 \$5467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44647 \$153 \$5031 \$5520 \$5338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44648 \$153 \$5901 \$4179 \$5742 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$44649 \$153 \$5592 \$5205 \$5564 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44651 \$153 \$5743 \$5519 \$5013 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44652 \$16 \$4229 \$16 \$153 \$5845 VNB sky130_fd_sc_hd__inv_1
X$44653 \$153 \$5468 \$5287 \$5013 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44656 \$153 \$5846 \$4616 \$5847 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$44657 \$153 \$5651 \$5669 \$5338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44658 \$16 \$4421 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44659 \$16 \$4178 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44660 \$153 \$5955 \$5390 \$5623 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44661 \$16 \$4178 \$16 \$153 \$5623 VNB sky130_fd_sc_hd__inv_1
X$44662 \$16 \$5338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44664 \$153 \$5848 \$5406 \$6032 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44665 \$153 \$5744 \$5069 \$5623 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44667 \$16 \$4421 \$5713 \$5827 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$44668 \$153 \$5745 \$5096 \$5623 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44669 \$153 \$5849 \$5388 \$5827 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$44670 \$153 \$5746 \$5519 \$5623 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44671 \$16 \$5772 \$16 \$153 \$5186 VNB sky130_fd_sc_hd__clkbuf_2
X$44673 \$153 \$5850 \$5653 \$5478 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44674 \$16 \$5772 \$16 \$153 \$5713 VNB sky130_fd_sc_hd__clkbuf_2
X$44675 \$153 \$5670 \$5209 \$5595 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44676 \$153 \$5594 \$5519 \$5170 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44677 \$16 \$5772 \$16 \$153 \$5900 VNB sky130_fd_sc_hd__clkbuf_2
X$44678 \$16 \$5478 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44679 \$153 \$5851 \$5653 \$5232 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44681 \$16 \$4421 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44683 \$153 \$5671 \$5096 \$5595 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44685 \$16 \$5232 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44686 \$153 \$5814 \$5653 \$5467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44687 \$153 \$5672 \$5287 \$5595 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44688 \$16 \$5765 \$16 \$153 \$3064 VNB sky130_fd_sc_hd__clkbuf_2
X$44689 \$16 \$5765 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44690 \$16 \$5467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44692 \$153 \$5445 \$5519 \$5283 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44694 \$153 \$5814 \$5406 \$5595 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44695 \$153 \$5725 \$5673 \$5338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44696 \$16 \$3064 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44697 \$153 \$5828 \$5406 \$5852 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44698 \$153 \$5829 \$5096 \$5852 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44699 \$16 \$4106 \$16 \$153 \$5726 VNB sky130_fd_sc_hd__inv_1
X$44701 \$16 \$5772 \$16 \$153 \$5479 VNB sky130_fd_sc_hd__clkbuf_2
X$44702 \$16 \$4106 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44703 \$16 \$4146 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44704 \$16 \$5338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44706 \$153 \$5853 \$5673 \$5467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44708 \$153 \$5654 \$5673 \$5324 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44709 \$16 \$5467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44710 \$153 \$5748 \$5205 \$5726 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44711 \$16 \$3886 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44714 \$153 \$5930 \$5390 \$5726 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44715 \$16 \$5324 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44716 \$16 \$3949 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44717 \$16 \$3658 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44720 \$153 \$5794 \$5549 \$5478 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44721 \$153 \$5854 \$5549 \$5469 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44723 \$153 \$5773 \$5549 \$5467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44725 \$153 \$5675 \$5205 \$5631 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44726 \$153 \$5773 \$5406 \$5631 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44727 \$153 \$5794 \$5390 \$5631 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44728 \$153 \$5539 \$5209 \$5631 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44729 \$16 \$5467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44730 \$16 \$4712 \$16 \$153 \$5815 VNB sky130_fd_sc_hd__inv_1
X$44731 \$16 \$4712 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44733 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44734 \$153 \$5855 \$5830 \$5232 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44735 \$153 \$5774 \$5519 \$5815 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44736 \$153 \$3343 \$1482 \$5755 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44737 \$16 \$5232 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44738 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$44739 \$153 \$5816 \$5830 \$5338 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44741 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44742 \$16 \$5500 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44743 \$16 \$5755 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44745 \$16 \$5795 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44746 \$16 \$5338 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44747 \$153 \$5816 \$5209 \$5815 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44748 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44749 \$153 \$3156 \$1482 \$5775 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44751 \$153 \$5749 \$5755 \$5471 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44753 \$153 \$5817 \$5632 \$5819 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44754 \$16 \$5796 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44756 \$153 \$5678 \$5625 \$5471 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44757 \$153 \$5879 \$5775 \$5471 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44758 \$153 \$5817 \$6200 \$5471 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44759 \$16 \$5775 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44760 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$44761 \$16 \$5819 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44763 \$153 \$153 \$5881 \$5568 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44764 \$153 \$153 \$5795 \$5568 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44767 \$153 \$5776 \$5632 \$5834 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44768 \$153 \$5933 \$5795 \$5471 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44769 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$44770 \$153 \$5776 \$5881 \$5471 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44771 \$16 \$5834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44775 \$16 \$5856 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44776 \$153 \$5750 \$5679 \$5796 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44777 \$153 \$5777 \$5679 \$5856 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44779 \$16 \$5819 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44780 \$16 \$3870 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44781 \$153 \$5857 \$5679 \$5819 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44782 \$16 \$4324 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44783 \$16 \$5714 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44785 \$153 \$5750 \$5775 \$5340 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44786 \$153 \$5777 \$5795 \$5340 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44787 \$153 \$5858 \$5679 \$5834 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44788 \$153 \$5751 \$5755 \$5340 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44789 \$16 \$5819 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44790 \$16 \$5714 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44792 \$16 \$3870 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44793 \$153 \$5779 \$5655 \$5819 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44795 \$153 \$5778 \$5795 \$5571 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44796 \$153 \$5779 \$6200 \$5571 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44798 \$16 \$5834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44799 \$153 \$5859 \$5655 \$5834 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44800 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$44803 \$153 \$5780 \$5775 \$5571 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44804 \$153 \$5780 \$5655 \$5796 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44805 \$153 \$5766 \$5470 \$5472 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44806 \$153 \$5766 \$5552 \$5702 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44807 \$16 \$5796 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44808 \$16 \$5702 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44811 \$153 \$5860 \$5552 \$5819 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44812 \$153 \$5752 \$5552 \$5796 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44813 \$153 \$5861 \$5552 \$5856 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44814 \$16 \$5796 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44815 \$16 \$3929 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44817 \$153 \$5752 \$5775 \$5472 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44818 \$16 \$5856 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44820 \$16 \$5856 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44821 \$153 \$5818 \$5633 \$5834 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44823 \$153 \$5797 \$5633 \$5856 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44824 \$16 \$5834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44825 \$153 \$5781 \$5775 \$5624 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44828 \$16 \$5819 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44829 \$153 \$5820 \$5633 \$5819 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44831 \$16 \$4011 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44832 \$16 \$4011 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44833 \$16 \$4011 \$16 \$153 \$5624 VNB sky130_fd_sc_hd__inv_1
X$44835 \$16 \$4258 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44836 \$153 \$5753 \$5755 \$5624 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44837 \$153 \$5820 \$6200 \$5624 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44842 \$153 \$5821 \$5656 \$5834 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44843 \$153 \$5798 \$5656 \$5856 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44844 \$153 \$5821 \$5881 \$5727 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44845 \$153 \$5682 \$5470 \$5727 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44847 \$16 \$5819 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44848 \$16 \$5906 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44849 \$16 \$4016 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44851 \$153 \$5862 \$5656 \$5819 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44852 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$44853 \$153 \$5754 \$5755 \$5727 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44855 \$16 \$5528 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44857 \$16 \$5819 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44858 \$153 \$5782 \$5658 \$5819 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44859 \$16 \$4152 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44860 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$44861 \$16 \$5356 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44862 \$16 \$5236 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44865 \$16 \$5799 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44866 \$16 \$5834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44867 \$153 \$5863 \$5658 \$5834 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44868 \$153 \$5782 \$6200 \$5434 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44869 \$16 \$4092 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44870 \$16 \$5906 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44871 \$16 \$5906 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44872 \$153 \$5783 \$5775 \$5434 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44874 \$16 \$3834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44875 \$16 \$5819 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44876 \$16 \$5702 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44879 \$16 \$5856 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44880 \$153 \$5756 \$5634 \$5856 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44881 \$153 \$5822 \$5634 \$5819 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44882 \$153 \$5756 \$5795 \$5574 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44883 \$153 \$5822 \$6200 \$5574 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44885 \$16 \$5194 \$5235 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$44887 \$153 \$5684 \$5625 \$5574 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44888 \$16 \$5194 \$5799 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$44890 \$153 \$5864 \$5634 \$5796 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44891 \$16 \$5194 \$5473 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$44893 \$16 \$4092 \$16 \$153 \$5574 VNB sky130_fd_sc_hd__inv_1
X$44895 \$153 \$5784 \$5755 \$5574 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44896 \$16 \$5796 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44897 \$16 \$4760 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44898 \$16 \$3983 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44899 \$16 \$5627 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44902 \$16 \$5484 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44904 \$153 \$153 \$5074 \$5715 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44905 \$16 \$16 \$153 VNB sky130_fd_sc_hd__conb_1
X$44906 \$153 \$153 \$5806 \$5715 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44907 \$153 \$153 \$5484 \$5715 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44908 \$153 \$153 \$5509 \$5715 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44909 \$153 \$153 \$5627 \$5715 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44910 \$16 \$5635 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44911 \$16 \$5480 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44913 \$16 \$5938 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44914 \$16 \$4324 \$16 \$153 \$5823 VNB sky130_fd_sc_hd__inv_1
X$44916 \$16 \$5887 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44918 \$16 \$5718 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44919 \$153 \$5757 \$5576 \$5887 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44920 \$153 \$5716 \$5576 \$5718 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44921 \$153 \$5962 \$5074 \$5823 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44922 \$16 \$5963 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44923 \$16 \$5541 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44924 \$16 \$5767 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44926 \$153 \$5785 \$5576 \$5767 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44927 \$153 \$5757 \$5627 \$5474 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44929 \$153 \$5785 \$5575 \$5474 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44931 \$16 \$5609 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44932 \$153 \$5506 \$5717 \$5609 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44933 \$16 \$5636 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44934 \$16 \$4126 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44935 \$16 \$4139 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44939 \$153 \$5758 \$5509 \$5475 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44941 \$16 \$5786 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44942 \$153 \$5800 \$5532 \$5786 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44943 \$16 \$5579 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44944 \$153 \$5865 \$5717 \$5579 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44945 \$153 \$5659 \$5509 \$5611 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44947 \$153 \$5800 \$5635 \$5611 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44948 \$16 \$5767 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44949 \$153 \$5801 \$5532 \$5767 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44951 \$153 \$5866 \$5532 \$5887 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44952 \$16 \$4560 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44953 \$153 \$5801 \$5575 \$5611 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44957 \$153 \$5759 \$5938 \$5614 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44959 \$153 \$5824 \$5835 \$5609 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44960 \$153 \$5802 \$5533 \$5767 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44962 \$16 \$4432 \$16 \$153 \$5867 VNB sky130_fd_sc_hd__inv_1
X$44963 \$16 \$5767 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44965 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$44966 \$153 \$5824 \$5074 \$5867 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44967 \$16 \$5786 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44968 \$153 \$5803 \$5533 \$5786 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44969 \$153 \$5802 \$5575 \$5614 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44971 \$153 \$5803 \$5635 \$5614 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44972 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$44974 \$16 \$5264 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44976 \$16 \$5718 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44977 \$16 \$5887 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44978 \$153 \$5868 \$5578 \$5718 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44979 \$153 \$5804 \$5578 \$5887 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44980 \$153 \$5804 \$5627 \$5559 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44982 \$16 \$5786 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44983 \$16 \$5767 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44984 \$153 \$5760 \$5578 \$5767 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44986 \$153 \$5825 \$5578 \$5786 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44987 \$153 \$5760 \$5575 \$5559 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44988 \$153 \$5825 \$5635 \$5559 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44990 \$16 \$3567 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44992 \$16 \$5767 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44993 \$16 \$5786 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44996 \$153 \$5831 \$5637 \$5767 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$44997 \$16 \$4016 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$44998 \$153 \$5761 \$5635 \$5511 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$44999 \$153 \$5831 \$5575 \$5511 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45000 \$16 \$5636 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45001 \$16 \$5887 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45002 \$16 \$5963 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45004 \$153 \$5805 \$5637 \$5963 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45005 \$16 \$3567 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45006 \$16 \$4092 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45007 \$16 \$5718 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45009 \$153 \$5787 \$5637 \$5718 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45010 \$153 \$5805 \$5806 \$5511 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45011 \$16 \$5579 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45012 \$153 \$5787 \$5938 \$5511 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45013 \$153 \$5788 \$5617 \$5579 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45015 \$153 \$5788 \$5484 \$5692 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45016 \$153 \$5789 \$5617 \$5963 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45017 \$153 \$5719 \$5617 \$5718 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45018 \$16 \$5963 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45019 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$45020 \$153 \$5789 \$5806 \$5692 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45023 \$16 \$5887 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45024 \$153 \$5583 \$5617 \$5887 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45025 \$153 \$5411 \$5617 \$5609 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45026 \$153 \$5869 \$5509 \$5692 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45027 \$16 \$5609 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45028 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$45030 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$45031 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$45032 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$45033 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$45034 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$45035 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$45036 \$153 \$1887 \$2009 \$1762 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45037 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$45039 \$153 \$1785 \$1873 \$1658 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45040 \$153 \$1786 \$1873 \$1687 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45041 \$16 \$1658 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45042 \$16 \$1687 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45045 \$153 \$1975 \$1943 \$1762 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45047 \$153 \$1836 \$1873 \$1795 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45048 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$45049 \$16 \$753 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45050 \$153 \$1873 \$531 \$1814 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$45051 \$153 \$1836 \$1815 \$1762 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45053 \$16 \$1795 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45055 \$16 \$264 \$16 \$153 \$1762 VNB sky130_fd_sc_hd__inv_1
X$45056 \$153 \$1791 \$1774 \$1687 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45057 \$16 \$1430 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45058 \$153 \$1977 \$1774 \$1980 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45059 \$16 \$1687 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45060 \$153 \$1837 \$1774 \$1795 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45061 \$16 \$1980 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45062 \$16 \$1480 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45064 \$153 \$1976 \$1792 \$1669 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45065 \$153 \$1838 \$1763 \$1687 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45067 \$16 \$582 \$16 \$153 \$1537 VNB sky130_fd_sc_hd__inv_1
X$45068 \$153 \$1790 \$1763 \$1658 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45069 \$16 \$263 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45072 \$153 \$1838 \$1792 \$1789 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45073 \$16 \$1687 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45074 \$16 \$1658 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45075 \$16 \$1686 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45076 \$16 \$1795 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45077 \$16 \$754 \$16 \$153 \$1789 VNB sky130_fd_sc_hd__inv_1
X$45078 \$153 \$1978 \$1888 \$1795 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45080 \$153 \$1839 \$1888 \$1687 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45081 \$16 \$279 \$16 \$153 \$1861 VNB sky130_fd_sc_hd__inv_1
X$45083 \$153 \$1837 \$1815 \$1537 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45084 \$153 \$1977 \$2009 \$1537 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45085 \$153 \$1978 \$1815 \$1861 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45086 \$153 \$1839 \$1792 \$1861 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45088 \$153 \$1889 \$1547 \$1861 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45089 \$153 \$1890 \$1963 \$1658 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45091 \$153 \$1794 \$1963 \$1687 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45092 \$16 \$1658 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45094 \$16 \$1168 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45095 \$153 \$1891 \$1963 \$1795 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45096 \$153 \$1890 \$1547 \$1793 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45098 \$153 \$1891 \$1815 \$1793 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45100 \$16 \$280 \$16 \$153 \$1793 VNB sky130_fd_sc_hd__inv_1
X$45101 \$16 \$1795 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45102 \$153 \$1892 \$1766 \$1658 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45103 \$16 \$1687 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45104 \$16 \$1576 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45106 \$153 \$1862 \$1766 \$1795 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45107 \$153 \$1979 \$1766 \$1980 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45110 \$153 \$1862 \$1815 \$1767 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45111 \$16 \$1658 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45112 \$153 \$1892 \$1547 \$1767 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45114 \$153 \$1893 \$1675 \$1795 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45115 \$153 \$1840 \$1675 \$1687 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45117 \$16 \$1942 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45119 \$153 \$1947 \$1675 \$1980 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45120 \$153 \$1893 \$1815 \$1796 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45121 \$153 \$1733 \$1547 \$1796 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45122 \$153 \$1947 \$2009 \$1796 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45123 \$16 \$356 \$16 \$153 \$1796 VNB sky130_fd_sc_hd__inv_1
X$45125 \$16 \$1980 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45126 \$153 \$1917 \$1676 \$1795 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45127 \$16 \$2006 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45128 \$153 \$1948 \$1676 \$2006 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45129 \$16 \$1795 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45130 \$16 \$356 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45132 \$16 \$1942 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45133 \$153 \$1748 \$1792 \$1670 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45134 \$16 \$1980 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45135 \$16 \$1522 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45136 \$16 \$899 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45138 \$153 \$1948 \$1943 \$1670 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45140 \$153 \$1691 \$1797 \$1795 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45141 \$153 \$1917 \$1815 \$1670 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45142 \$153 \$1749 \$1792 \$1671 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45143 \$16 \$1795 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45144 \$16 \$351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45145 \$16 \$1551 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45146 \$16 \$2006 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45147 \$153 \$1949 \$1797 \$2006 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45149 \$153 \$1841 \$1797 \$1658 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45150 \$153 \$1949 \$1943 \$1671 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45151 \$153 \$1841 \$1547 \$1671 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45152 \$16 \$1658 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45153 \$16 \$2647 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45154 \$16 \$351 \$16 \$153 \$1671 VNB sky130_fd_sc_hd__inv_1
X$45156 \$16 \$1775 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45159 \$16 \$351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45160 \$16 \$584 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45161 \$153 \$1798 \$1768 \$1816 \$1799 \$1777 \$16 \$16 VNB
+ sky130_fd_sc_hd__nor4b_2
X$45162 \$153 \$1776 \$1799 \$1777 \$1816 \$1768 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$45163 \$153 \$1816 \$1799 \$1964 \$1768 \$1777 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$45164 \$153 \$1768 \$1799 \$1800 \$1816 \$1777 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$45165 \$16 \$1964 \$16 \$153 \$710 VNB sky130_fd_sc_hd__clkbuf_2
X$45167 \$16 \$1918 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45168 \$16 \$1981 \$16 \$153 \$1013 VNB sky130_fd_sc_hd__clkbuf_2
X$45171 \$16 \$1874 \$16 \$153 \$380 VNB sky130_fd_sc_hd__clkbuf_2
X$45172 \$16 \$1894 \$16 \$153 \$279 VNB sky130_fd_sc_hd__clkbuf_2
X$45173 \$153 \$1894 \$1875 \$1842 \$1863 \$2038 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$45174 \$153 \$1874 \$1863 \$1875 \$2038 \$1842 \$16 \$16 VNB
+ sky130_fd_sc_hd__nor4b_2
X$45175 \$153 \$1504 \$1595 \$1660 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$45176 \$153 \$1875 \$1863 \$1801 \$2038 \$1842 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$45179 \$153 \$1919 \$454 \$1817 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$45180 \$153 \$2039 \$531 \$1982 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$45181 \$16 \$1595 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45182 \$16 \$264 \$16 \$153 \$1944 VNB sky130_fd_sc_hd__inv_1
X$45183 \$16 \$59 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45185 \$153 \$1865 \$1895 \$1864 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45186 \$153 \$1950 \$1919 \$1965 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45188 \$153 \$1865 \$1919 \$1923 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45189 \$153 \$1950 \$1806 \$1864 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45190 \$153 \$1983 \$1924 \$1864 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45192 \$153 \$1920 \$1919 \$1805 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45193 \$16 \$1965 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45194 \$16 \$264 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45196 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$45197 \$153 \$1984 \$1471 \$1944 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45198 \$16 \$1805 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45199 \$153 \$1661 \$347 \$1633 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45200 \$153 \$1803 \$1779 \$2042 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45201 \$153 \$1920 \$1703 \$1864 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45203 \$16 \$979 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45205 \$16 \$754 \$16 \$153 \$1483 VNB sky130_fd_sc_hd__inv_1
X$45206 \$16 \$2042 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45208 \$16 \$1923 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45209 \$153 \$1507 \$1779 \$1845 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45211 \$153 \$1769 \$1779 \$1965 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45213 \$153 \$1921 \$541 \$1896 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$45214 \$16 \$1965 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45215 \$16 \$1845 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45216 \$16 \$1966 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45218 \$16 \$279 \$1966 \$1896 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$45219 \$153 \$1554 \$1921 \$1923 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45220 \$153 \$1951 \$1921 \$1965 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45221 \$16 \$279 \$16 \$153 \$1922 VNB sky130_fd_sc_hd__inv_1
X$45222 \$153 \$1951 \$1806 \$1922 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45223 \$16 \$710 \$16 \$153 \$1866 VNB sky130_fd_sc_hd__inv_1
X$45225 \$153 \$1698 \$1697 \$1923 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45226 \$153 \$2013 \$1703 \$1922 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45228 \$153 \$1985 \$1697 \$1965 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45229 \$153 \$1818 \$1703 \$1866 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45230 \$153 \$1819 \$1471 \$1866 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45232 \$16 \$1965 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45233 \$16 \$2042 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45236 \$153 \$1945 \$1820 \$1965 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45237 \$153 \$1843 \$1820 \$1845 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45238 \$153 \$1952 \$1820 \$1923 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45239 \$16 \$323 \$16 \$153 \$1844 VNB sky130_fd_sc_hd__inv_1
X$45240 \$16 \$1845 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45242 \$153 \$1945 \$1806 \$1844 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45243 \$153 \$1821 \$1703 \$1844 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45244 \$16 \$1805 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45245 \$16 \$1923 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45246 \$16 \$1845 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45248 \$153 \$1702 \$1700 \$1805 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45249 \$153 \$1952 \$1895 \$1844 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45252 \$16 \$1923 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45254 \$153 \$1897 \$1700 \$1965 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45255 \$153 \$1867 \$1924 \$1822 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45256 \$16 \$1805 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45257 \$16 \$1845 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45258 \$153 \$1897 \$1806 \$1822 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45259 \$16 \$380 \$1966 \$1823 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$45261 \$16 \$1965 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45262 \$153 \$1953 \$1770 \$1965 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45264 \$16 \$684 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45265 \$16 \$380 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45266 \$153 \$1780 \$505 \$1824 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$45267 \$153 \$1807 \$1895 \$1822 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45269 \$16 \$1845 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45270 \$153 \$1846 \$1770 \$1845 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45271 \$16 \$1965 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45272 \$16 \$1966 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45273 \$16 \$1966 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45275 \$153 \$1986 \$1954 \$1752 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45276 \$153 \$1754 \$1703 \$1752 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45277 \$153 \$1953 \$1806 \$1752 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45278 \$153 \$1753 \$1895 \$1752 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45279 \$153 \$1987 \$1954 \$1704 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45281 \$16 \$351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45283 \$153 \$1847 \$1780 \$1965 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45284 \$16 \$1508 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45285 \$16 \$1508 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45286 \$153 \$1898 \$1780 \$1805 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45287 \$153 \$1847 \$1806 \$1704 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45288 \$16 \$1805 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45289 \$16 \$2199 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45290 \$153 \$1898 \$1703 \$1704 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45291 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$45293 \$153 \$1988 \$1967 \$1805 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45295 \$16 \$54 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45296 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45297 \$153 \$1925 \$1482 \$389 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45298 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45299 \$153 \$1989 \$1482 \$54 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45302 \$153 \$1755 \$1471 \$1704 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45303 \$153 \$1990 \$1967 \$1965 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45304 \$16 \$1965 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45305 \$16 \$389 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45306 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$45307 \$153 \$1642 \$1876 \$1969 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45308 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$45309 \$16 \$253 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45312 \$153 \$1557 \$1876 \$1879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45313 \$153 \$2245 \$1482 \$388 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45314 \$16 \$1879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45315 \$153 \$1955 \$1876 \$1878 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45316 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45317 \$16 \$1969 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45318 \$16 \$388 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45321 \$153 \$1848 \$1876 \$1756 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45322 \$153 \$1876 \$387 \$1877 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$45323 \$16 \$426 \$1968 \$1877 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$45324 \$16 \$1878 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45325 \$16 \$1878 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45326 \$16 \$2105 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45327 \$153 \$1849 \$1781 \$1878 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45328 \$16 \$266 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45329 \$16 \$1756 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45331 \$153 \$1808 \$1781 \$1756 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45332 \$153 \$1849 \$1868 \$1679 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45333 \$16 \$2016 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45334 \$153 \$1899 \$1781 \$1879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45335 \$16 \$1879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45337 \$16 \$265 \$1929 \$1926 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$45340 \$16 \$399 \$16 \$153 \$1679 VNB sky130_fd_sc_hd__inv_1
X$45341 \$153 \$1899 \$1558 \$1679 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45342 \$153 \$1781 \$595 \$1740 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$45343 \$16 \$424 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45344 \$153 \$1900 \$423 \$1926 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$45346 \$16 \$1878 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45347 \$16 \$964 \$1968 \$1946 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$45349 \$153 \$1901 \$1900 \$1878 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45350 \$153 \$1850 \$1900 \$1756 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45351 \$16 \$2105 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45352 \$153 \$1901 \$1868 \$1771 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45353 \$16 \$1969 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45354 \$153 \$1828 \$1900 \$1969 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45355 \$16 \$1879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45357 \$153 \$1809 \$1900 \$1879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45358 \$16 \$265 \$16 \$153 \$1771 VNB sky130_fd_sc_hd__inv_1
X$45360 \$16 \$798 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45361 \$153 \$1880 \$856 \$1927 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$45362 \$16 \$798 \$1968 \$1927 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$45363 \$16 \$1878 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45364 \$153 \$1851 \$1880 \$1878 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45366 \$153 \$1709 \$1880 \$1756 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45367 \$153 \$1851 \$1868 \$1674 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45368 \$153 \$1991 \$1880 \$1879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45369 \$16 \$1879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45370 \$16 \$423 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45371 \$16 \$399 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45372 \$16 \$1760 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45375 \$153 \$1928 \$591 \$1902 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$45376 \$153 \$1810 \$1880 \$1969 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45377 \$153 \$1562 \$1928 \$1879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45378 \$16 \$151 \$1929 \$1902 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$45379 \$16 \$1929 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45382 \$16 \$151 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45383 \$16 \$1514 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45384 \$16 \$1879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45385 \$16 \$1585 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45387 \$16 \$1446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45388 \$16 \$1756 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45389 \$153 \$1254 \$1627 \$1829 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$45390 \$153 \$1713 \$1928 \$1756 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45391 \$16 \$424 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45392 \$16 \$1929 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45393 \$153 \$1992 \$1993 \$1542 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45394 \$16 \$1879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45396 \$16 \$306 \$1929 \$1830 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$45398 \$16 \$1878 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45399 \$153 \$1852 \$1903 \$1879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45400 \$153 \$1994 \$1903 \$1878 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45401 \$153 \$1853 \$1903 \$1756 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45402 \$16 \$1756 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45404 \$16 \$1969 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45406 \$153 \$1904 \$1903 \$1969 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45407 \$153 \$1853 \$1712 \$1759 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45408 \$16 \$1969 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45409 \$153 \$1904 \$1613 \$1759 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45410 \$153 \$1995 \$1854 \$1969 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45412 \$153 \$1930 \$1854 \$1878 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45413 \$16 \$1878 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45414 \$153 \$1930 \$1868 \$1996 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45415 \$153 \$1931 \$1854 \$1756 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45416 \$16 \$1756 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45417 \$153 \$1932 \$1558 \$1996 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45419 \$153 \$1931 \$1712 \$1996 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45420 \$153 \$1932 \$1854 \$1879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45421 \$153 \$1881 \$1970 \$1782 \$1831 \$1812 \$16 \$16 VNB
+ sky130_fd_sc_hd__nor4b_2
X$45422 \$16 \$1881 \$16 \$153 \$829 VNB sky130_fd_sc_hd__clkbuf_2
X$45423 \$153 \$1782 \$1970 \$1884 \$1831 \$1812 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$45424 \$16 \$1882 \$16 \$153 \$265 VNB sky130_fd_sc_hd__clkbuf_2
X$45426 \$16 \$724 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45428 \$16 \$1593 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45429 \$16 \$1869 \$16 \$153 \$1044 VNB sky130_fd_sc_hd__clkbuf_2
X$45430 \$16 \$1997 \$16 \$153 \$426 VNB sky130_fd_sc_hd__clkbuf_2
X$45431 \$153 \$1869 \$1971 \$1855 \$1883 \$1905 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$45432 \$153 \$1997 \$1905 \$1883 \$1971 \$1855 \$16 \$16 VNB
+ sky130_fd_sc_hd__nor4b_2
X$45433 \$16 \$1884 \$16 \$153 \$306 VNB sky130_fd_sc_hd__clkbuf_2
X$45435 \$16 \$426 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45437 \$16 \$1933 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45438 \$16 \$426 \$1972 \$1956 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$45439 \$16 \$1601 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45440 \$16 \$371 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45441 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45443 \$153 \$1906 \$387 \$1956 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$45444 \$153 \$2774 \$1482 \$371 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45445 \$16 \$426 \$16 \$153 \$1999 VNB sky130_fd_sc_hd__inv_1
X$45447 \$16 \$1832 \$1933 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$45448 \$16 \$1832 \$1628 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$45449 \$16 \$1832 \$1647 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$45450 \$16 \$1832 \$1649 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$45451 \$153 \$1998 \$1906 \$1973 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45452 \$16 \$1832 \$1760 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$45454 \$16 \$2031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45455 \$16 \$964 \$1972 \$1856 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$45456 \$16 \$1784 \$116 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$45457 \$16 \$1784 \$998 \$153 \$16 VNB sky130_fd_sc_hd__clkbuf_1
X$45459 \$153 \$1957 \$1906 \$1960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45461 \$153 \$1934 \$1906 \$1860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45463 \$153 \$1957 \$2086 \$1999 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45464 \$16 \$399 \$1885 \$1907 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$45465 \$153 \$1935 \$595 \$1907 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$45466 \$153 \$1934 \$2000 \$1999 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45467 \$16 \$446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45468 \$16 \$178 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45469 \$153 \$1958 \$1974 \$1860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45470 \$16 \$265 \$1885 \$1908 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$45473 \$153 \$1909 \$423 \$1908 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$45474 \$153 \$1958 \$2000 \$2129 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45475 \$16 \$509 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45476 \$16 \$1885 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45477 \$16 \$1960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45478 \$153 \$1857 \$371 \$1651 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45480 \$16 \$1860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45481 \$153 \$1858 \$1909 \$1860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45483 \$16 \$265 \$16 \$153 \$1870 VNB sky130_fd_sc_hd__inv_1
X$45485 \$16 \$1973 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45486 \$153 \$1911 \$1909 \$1973 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45487 \$153 \$1910 \$2086 \$1870 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45488 \$153 \$1858 \$2000 \$1870 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45489 \$16 \$798 \$1972 \$2019 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$45491 \$16 \$1860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45492 \$153 \$1911 \$2056 \$1870 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45493 \$153 \$1959 \$2058 \$1860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45494 \$16 \$1972 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45495 \$153 \$1912 \$2056 \$2172 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45496 \$153 \$1959 \$2000 \$2172 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45497 \$153 \$1342 \$1708 \$1833 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$45498 \$16 \$1960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45500 \$153 \$2001 \$2058 \$1960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45501 \$16 \$354 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45503 \$153 \$1871 \$1936 \$2172 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45504 \$153 \$1886 \$591 \$1937 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$45505 \$16 \$151 \$1885 \$1937 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$45506 \$16 \$1514 \$1601 \$1859 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$45509 \$153 \$1834 \$371 \$1343 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45510 \$16 \$1960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45511 \$153 \$2002 \$1886 \$1960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45512 \$153 \$1938 \$608 \$1913 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$45513 \$16 \$306 \$1885 \$1913 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$45514 \$16 \$1973 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45516 \$16 \$1860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45517 \$153 \$1939 \$1886 \$1973 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45519 \$153 \$2003 \$1886 \$1860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45520 \$153 \$1492 \$1649 \$1914 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$45521 \$16 \$1599 \$1601 \$1914 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$45522 \$153 \$1961 \$2004 \$1973 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45525 \$16 \$829 \$16 \$153 \$1940 VNB sky130_fd_sc_hd__inv_1
X$45526 \$16 \$1973 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45527 \$16 \$829 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45528 \$16 \$1860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45529 \$153 \$1961 \$2056 \$1940 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45530 \$153 \$1746 \$371 \$1344 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45532 \$153 \$1941 \$2000 \$1940 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45533 \$153 \$1941 \$2004 \$1860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45535 \$16 \$1599 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45537 \$16 \$306 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45538 \$153 \$2005 \$2086 \$1940 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45539 \$153 \$1416 \$1627 \$1835 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$45540 \$16 \$306 \$16 \$153 \$1872 VNB sky130_fd_sc_hd__inv_1
X$45541 \$153 \$1915 \$1938 \$1860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45542 \$16 \$1860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45543 \$16 \$1627 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45544 \$16 \$1758 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45548 \$153 \$1915 \$2000 \$1872 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45549 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$45551 \$16 \$1960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45552 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$45553 \$153 \$1962 \$1938 \$1960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45554 \$16 \$446 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45555 \$153 \$1813 \$1416 \$446 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45557 \$153 \$1962 \$2086 \$1872 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45558 \$153 \$1916 \$1936 \$1872 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45559 \$153 \$2022 \$2056 \$1872 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45560 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$45561 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$45563 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$45564 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$45565 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$45566 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$45567 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$45568 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$45569 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$45571 \$153 \$4767 \$4469 \$3766 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45572 \$153 \$4629 \$4469 \$3709 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45573 \$16 \$3766 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45574 \$16 \$3709 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45575 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$45576 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$45577 \$153 \$4741 \$4469 \$3385 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45579 \$153 \$4767 \$3478 \$4372 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45580 \$16 \$4742 \$16 \$153 \$4372 VNB sky130_fd_sc_hd__inv_1
X$45581 \$153 \$4741 \$3394 \$4372 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45582 \$16 \$3385 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45583 \$16 \$4742 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45584 \$153 \$4576 \$3540 \$4372 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45585 \$153 \$4809 \$3540 \$4859 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45587 \$16 \$4902 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45589 \$153 \$4649 \$3422 \$4372 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45590 \$153 \$4768 \$4788 \$3709 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45591 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$45592 \$16 \$4579 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45593 \$153 \$4703 \$3307 \$4692 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45594 \$153 \$4768 \$3606 \$4692 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45596 \$16 \$3615 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45598 \$153 \$4810 \$4788 \$3474 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45599 \$153 \$4650 \$3307 \$4489 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45600 \$153 \$4704 \$3540 \$4692 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45601 \$16 \$3474 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45602 \$153 \$4705 \$4706 \$4579 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45603 \$16 \$4538 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45605 \$16 \$5080 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45606 \$153 \$4769 \$4614 \$3709 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45608 \$153 \$4652 \$4614 \$3615 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45609 \$153 \$4769 \$3606 \$4707 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45610 \$153 \$4651 \$3490 \$4707 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45611 \$16 \$3615 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45612 \$16 \$3473 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45613 \$16 \$3709 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45614 \$153 \$4653 \$3540 \$4707 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45615 \$16 \$4479 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45617 \$153 \$4546 \$4789 \$3615 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45618 \$153 \$4652 \$3307 \$4707 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45619 \$153 \$4708 \$3490 \$4693 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45621 \$153 \$4811 \$4617 \$3615 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45622 \$16 \$3615 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45625 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$45627 \$16 \$3615 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45628 \$16 \$3616 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45629 \$153 \$4595 \$3394 \$4527 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45630 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$45631 \$16 \$4812 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45632 \$153 \$4813 \$4865 \$3615 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45633 \$153 \$4617 \$4812 \$4654 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$45635 \$153 \$4770 \$4617 \$3571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45636 \$153 \$4655 \$4617 \$3709 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45637 \$153 \$4770 \$3422 \$4527 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45638 \$153 \$4655 \$3606 \$4527 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45639 \$16 \$4621 \$16 \$153 \$4527 VNB sky130_fd_sc_hd__inv_1
X$45643 \$153 \$4630 \$4386 \$3385 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45644 \$153 \$4743 \$4386 \$3571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45645 \$153 \$4743 \$3422 \$4373 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45646 \$153 \$4388 \$4867 \$3615 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45647 \$16 \$3571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45650 \$16 \$3385 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45652 \$16 \$4600 \$16 \$153 \$4373 VNB sky130_fd_sc_hd__inv_1
X$45653 \$153 \$4386 \$5230 \$4657 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$45655 \$153 \$4656 \$3307 \$4373 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45656 \$16 \$3615 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45658 \$153 \$4709 \$3389 \$4359 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45659 \$153 \$4790 \$3490 \$4359 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45661 \$153 \$4786 \$3540 \$4359 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45662 \$153 \$4744 \$4390 \$3385 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45664 \$16 \$3474 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45665 \$153 \$4814 \$4791 \$3474 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45666 \$153 \$4658 \$3490 \$4329 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45667 \$153 \$4710 \$4390 \$3571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45669 \$153 \$4744 \$3394 \$4329 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45671 \$153 \$4390 \$5065 \$4745 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$45672 \$153 \$4710 \$3422 \$4329 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45673 \$16 \$4712 \$4012 \$4745 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$45674 \$153 \$4713 \$4711 \$3473 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45677 \$16 \$3474 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45678 \$153 \$4746 \$4711 \$3615 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45679 \$153 \$4771 \$4711 \$3474 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45680 \$153 \$4713 \$3540 \$4694 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45681 \$16 \$3615 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45683 \$16 \$4494 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45684 \$153 \$4771 \$3490 \$4694 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45685 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$45686 \$16 \$4792 \$16 \$153 \$3886 VNB sky130_fd_sc_hd__clkbuf_2
X$45688 \$16 \$4272 \$16 \$153 \$4659 VNB sky130_fd_sc_hd__clkbuf_2
X$45689 \$153 \$4792 \$4715 \$4659 \$4714 \$4598 \$16 \$16 VNB
+ sky130_fd_sc_hd__nor4b_2
X$45690 \$153 \$4659 \$4715 \$4747 \$4714 \$4598 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$45691 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$45692 \$16 \$4184 \$16 \$153 \$4715 VNB sky130_fd_sc_hd__clkbuf_2
X$45694 \$16 \$4660 \$16 \$153 \$4479 VNB sky130_fd_sc_hd__clkbuf_2
X$45696 \$16 \$4078 \$16 \$153 \$4661 VNB sky130_fd_sc_hd__clkbuf_2
X$45698 \$16 \$4184 \$16 \$153 \$4716 VNB sky130_fd_sc_hd__clkbuf_2
X$45700 \$16 \$4793 \$16 \$153 \$4320 VNB sky130_fd_sc_hd__clkbuf_2
X$45701 \$16 \$4272 \$16 \$153 \$4717 VNB sky130_fd_sc_hd__clkbuf_2
X$45702 \$153 \$4794 \$4716 \$4662 \$4717 \$4661 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$45703 \$153 \$4716 \$4661 \$4748 \$4717 \$4662 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$45704 \$153 \$4540 \$4812 \$4718 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$45705 \$16 \$4794 \$16 \$153 \$4742 VNB sky130_fd_sc_hd__clkbuf_2
X$45706 \$16 \$4275 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45708 \$16 \$4621 \$4275 \$4718 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$45710 \$153 \$4815 \$4599 \$3621 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45711 \$153 \$4749 \$4599 \$3572 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45712 \$16 \$4902 \$16 \$153 \$4529 VNB sky130_fd_sc_hd__inv_1
X$45713 \$16 \$3572 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45714 \$16 \$3621 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45715 \$16 \$3572 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45717 \$153 \$4772 \$4599 \$3543 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45718 \$153 \$4750 \$4599 \$3573 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45719 \$153 \$4772 \$3556 \$4529 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45720 \$153 \$4663 \$3101 \$4633 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45721 \$16 \$3543 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45722 \$16 \$3573 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45725 \$153 \$4719 \$4599 \$3620 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45727 \$153 \$4816 \$4599 \$3492 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45728 \$153 \$4719 \$3645 \$4529 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45729 \$153 \$4584 \$3435 \$4529 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45730 \$16 \$3620 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45731 \$16 \$3492 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45734 \$153 \$4664 \$3435 \$4633 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45736 \$153 \$4695 \$4540 \$3543 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45738 \$153 \$4795 \$3079 \$4796 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45739 \$153 \$4695 \$3556 \$4633 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45740 \$153 \$4787 \$3354 \$4796 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45741 \$16 \$3543 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45743 \$153 \$4787 \$4873 \$3492 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45744 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$45745 \$153 \$4553 \$4398 \$3492 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45746 \$16 \$3492 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45747 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$45748 \$16 \$3492 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45749 \$153 \$4773 \$4797 \$3573 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45750 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$45751 \$16 \$3480 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45753 \$153 \$4555 \$4398 \$3543 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45754 \$153 \$4817 \$3435 \$4818 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45755 \$16 \$3543 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45757 \$153 \$4773 \$3079 \$4818 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45758 \$16 \$3386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45759 \$153 \$4665 \$4622 \$3386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45763 \$153 \$4819 \$3608 \$4818 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45764 \$153 \$4603 \$3608 \$4530 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45765 \$16 \$3620 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45766 \$153 \$4774 \$4622 \$3543 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45767 \$153 \$4665 \$3435 \$4530 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45770 \$153 \$4774 \$3556 \$4530 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45771 \$153 \$4604 \$3645 \$4530 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45772 \$16 \$3620 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45773 \$153 \$4541 \$5230 \$4666 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$45774 \$16 \$5230 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45776 \$153 \$4820 \$3079 \$4798 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45777 \$153 \$4751 \$4541 \$3386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45778 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$45780 \$153 \$4821 \$4875 \$3492 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45781 \$153 \$4667 \$3645 \$4498 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45782 \$153 \$4751 \$3435 \$4498 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45783 \$16 \$3386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45784 \$16 \$3492 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45786 \$16 \$4668 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45787 \$153 \$4775 \$4541 \$3480 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45789 \$153 \$4670 \$4541 \$3572 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45790 \$153 \$4586 \$3556 \$4498 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45791 \$153 \$4670 \$3101 \$4498 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45792 \$16 \$3480 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45793 \$16 \$3492 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45794 \$16 \$3572 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45795 \$16 \$4822 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45796 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$45798 \$153 \$4720 \$4876 \$3386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45799 \$153 \$4402 \$4480 \$3386 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45800 \$153 \$4823 \$3608 \$4696 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45801 \$153 \$4720 \$3435 \$4696 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45802 \$16 \$3386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45804 \$16 \$3386 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45805 \$153 \$4752 \$4480 \$3543 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45806 \$153 \$4404 \$5228 \$4824 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$45807 \$153 \$4752 \$3556 \$4363 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45808 \$16 \$3543 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45809 \$16 \$3573 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45810 \$153 \$4671 \$4721 \$3573 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45812 \$16 \$4712 \$16 \$153 \$4776 VNB sky130_fd_sc_hd__inv_1
X$45815 \$153 \$4825 \$3645 \$5066 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45816 \$153 \$4671 \$3079 \$4776 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45817 \$153 \$4848 \$3504 \$4776 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45819 \$153 \$4672 \$3608 \$4501 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45820 \$153 \$4826 \$4721 \$3492 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45823 \$16 \$4869 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45824 \$153 \$4634 \$4721 \$3620 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45825 \$16 \$3572 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45826 \$153 \$4777 \$4721 \$3572 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45827 \$153 \$4635 \$4721 \$3543 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45828 \$16 \$3620 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45831 \$153 \$4777 \$3101 \$4776 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45832 \$16 \$3241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45833 \$16 \$3543 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45836 \$153 \$4778 \$4799 \$3731 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45837 \$153 \$4559 \$4481 \$3731 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45838 \$153 \$4800 \$3962 \$4801 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45840 \$16 \$3731 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45841 \$16 \$3731 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45842 \$153 \$4673 \$4481 \$3792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45843 \$153 \$4778 \$3788 \$4801 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45844 \$16 \$4780 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45845 \$153 \$4753 \$3919 \$4531 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45846 \$153 \$4753 \$4481 \$3791 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45848 \$16 \$4780 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45849 \$153 \$4802 \$3651 \$4801 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45850 \$16 \$4780 \$16 \$153 \$4531 VNB sky130_fd_sc_hd__inv_1
X$45852 \$153 \$4754 \$4722 \$3960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45853 \$16 \$4780 \$4166 \$4674 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$45855 \$153 \$4723 \$4722 \$3791 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45857 \$16 \$3960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45858 \$16 \$3814 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45859 \$153 \$4723 \$3919 \$4697 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45861 \$16 \$4759 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45862 \$16 \$3731 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45863 \$16 \$4048 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45864 \$153 \$4779 \$4722 \$3731 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45865 \$16 \$3852 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45866 \$153 \$4676 \$4722 \$3852 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45868 \$153 \$4779 \$3788 \$4697 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45869 \$153 \$4676 \$3763 \$4697 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45870 \$16 \$3960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45872 \$153 \$4755 \$4698 \$3852 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45873 \$153 \$4636 \$4698 \$3731 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45875 \$16 \$4560 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45876 \$153 \$4755 \$3763 \$4637 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45878 \$16 \$3814 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45879 \$16 \$4048 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45880 \$153 \$4757 \$4698 \$3814 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45881 \$153 \$4852 \$3716 \$4637 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45883 \$153 \$4677 \$3858 \$4637 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45884 \$16 \$4756 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45886 \$16 \$3731 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45888 \$16 \$4949 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45889 \$16 \$3814 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45890 \$16 \$3791 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45891 \$153 \$4623 \$4638 \$3731 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45892 \$153 \$4827 \$4638 \$3791 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45893 \$153 \$4757 \$3651 \$4637 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45894 \$153 \$4853 \$3763 \$4587 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45897 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$45898 \$16 \$3889 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45899 \$153 \$4758 \$4638 \$3889 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45901 \$16 \$4781 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45902 \$153 \$4678 \$3858 \$4587 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45903 \$153 \$4827 \$3919 \$4587 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45904 \$16 \$4475 \$16 \$153 \$4724 VNB sky130_fd_sc_hd__clkbuf_2
X$45905 \$153 \$4257 \$4609 \$4725 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$45906 \$16 \$4724 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45908 \$153 \$4758 \$3962 \$4587 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45910 \$16 \$4048 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45911 \$16 \$3791 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45912 \$153 \$4727 \$4726 \$4048 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45913 \$153 \$4679 \$4726 \$3791 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45914 \$153 \$4727 \$3858 \$4639 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45916 \$16 \$3792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45917 \$153 \$4640 \$4726 \$3814 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45918 \$16 \$3814 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45919 \$16 \$3731 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45920 \$153 \$4726 \$4803 \$4828 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$45921 \$153 \$4728 \$4726 \$3852 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45922 \$16 \$3960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45924 \$153 \$4829 \$4726 \$3731 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45925 \$16 \$3731 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45927 \$16 \$3792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45928 \$153 \$4699 \$4565 \$3792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45929 \$16 \$4803 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45931 \$16 \$4782 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45932 \$16 \$3792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45933 \$153 \$4783 \$4804 \$3792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45935 \$16 \$5158 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45936 \$16 \$4954 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45937 \$153 \$4680 \$3716 \$4532 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45938 \$153 \$4829 \$3788 \$4639 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45939 \$153 \$4699 \$3939 \$4532 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45940 \$16 \$3731 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45941 \$16 \$3567 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45942 \$16 \$4830 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45943 \$16 \$4830 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45944 \$153 \$4681 \$3763 \$4532 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45945 \$16 \$4831 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45947 \$16 \$4724 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45948 \$16 \$4724 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45949 \$16 \$4567 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45950 \$16 \$3814 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45951 \$16 \$3791 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45952 \$153 \$4682 \$3858 \$4532 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45953 \$153 \$4832 \$4804 \$3791 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45954 \$153 \$4729 \$3788 \$4700 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45955 \$16 \$4784 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45956 \$16 \$4567 \$16 \$153 \$4532 VNB sky130_fd_sc_hd__inv_1
X$45957 \$153 \$4684 \$3651 \$4532 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45959 \$153 \$4683 \$3919 \$4532 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45960 \$16 \$3814 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45961 \$16 \$2387 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45962 \$16 \$4805 \$16 \$153 \$4780 VNB sky130_fd_sc_hd__clkbuf_2
X$45963 \$16 \$4701 \$16 \$153 \$4093 VNB sky130_fd_sc_hd__clkbuf_2
X$45964 \$16 \$4347 \$16 \$153 \$4833 VNB sky130_fd_sc_hd__clkbuf_2
X$45965 \$16 \$4347 \$16 \$153 \$4641 VNB sky130_fd_sc_hd__clkbuf_2
X$45967 \$16 \$4834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45968 \$153 \$4685 \$4730 \$4610 \$4686 \$4641 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$45969 \$16 \$4589 \$16 \$153 \$4935 VNB sky130_fd_sc_hd__clkbuf_2
X$45970 \$16 \$4317 \$16 \$153 \$4730 VNB sky130_fd_sc_hd__clkbuf_2
X$45972 \$153 \$4701 \$4686 \$4610 \$4730 \$4641 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$45973 \$153 \$4805 \$4641 \$4610 \$4686 \$4730 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$45974 \$153 \$4686 \$4730 \$4533 \$4641 \$4610 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$45975 \$153 \$4730 \$4641 \$4732 \$4686 \$4610 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$45976 \$16 \$4610 \$4641 \$4686 \$4730 \$16 \$153 \$4534 VNB
+ sky130_fd_sc_hd__and4_2
X$45977 \$153 \$4686 \$4641 \$4835 \$4730 \$4610 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$45979 \$16 \$4759 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45980 \$16 \$3826 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45983 \$153 \$4611 \$4414 \$4643 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45984 \$153 \$4687 \$4731 \$3898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45985 \$153 \$4806 \$3860 \$4807 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45986 \$16 \$4732 \$16 \$153 \$4139 VNB sky130_fd_sc_hd__clkbuf_2
X$45987 \$16 \$4835 \$16 \$153 \$4415 VNB sky130_fd_sc_hd__clkbuf_2
X$45989 \$153 \$4688 \$4731 \$3691 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45990 \$16 \$3898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45993 \$153 \$4644 \$4731 \$3680 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$45994 \$153 \$4688 \$3142 \$4643 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$45995 \$16 \$3680 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45997 \$16 \$4129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45998 \$16 \$3691 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$45999 \$153 \$4645 \$4731 \$4129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46000 \$16 \$4760 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46002 \$16 \$3826 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46004 \$153 \$4733 \$4731 \$3826 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46005 \$153 \$4733 \$3893 \$4643 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46006 \$16 \$3898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46007 \$16 \$3721 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46008 \$153 \$4465 \$3860 \$4378 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46009 \$153 \$4761 \$4626 \$3721 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46012 \$16 \$3602 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46013 \$16 \$3680 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46014 \$153 \$4761 \$3676 \$4484 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46015 \$16 \$3064 \$16 \$153 \$4613 VNB sky130_fd_sc_hd__clkbuf_2
X$46016 \$153 \$4734 \$4626 \$3602 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46017 \$16 \$3064 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46018 \$153 \$4735 \$4626 \$3680 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46021 \$153 \$4735 \$3719 \$4484 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46022 \$153 \$4734 \$3565 \$4484 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46023 \$153 \$4689 \$4627 \$4129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46024 \$16 \$4057 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46025 \$16 \$4560 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46026 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$46027 \$153 \$4762 \$3142 \$4808 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46028 \$153 \$4762 \$4627 \$3691 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46031 \$16 \$3826 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46032 \$153 \$4785 \$4627 \$3826 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46033 \$153 \$4689 \$3986 \$4808 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46034 \$153 \$4785 \$3893 \$4808 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46036 \$16 \$4613 \$16 \$153 \$4736 VNB sky130_fd_sc_hd__clkbuf_2
X$46038 \$153 \$4690 \$4414 \$4808 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46040 \$16 \$4562 \$4736 \$4691 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$46042 \$153 \$4410 \$4737 \$3898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46043 \$16 \$3898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46044 \$16 \$3602 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46045 \$153 \$4642 \$4737 \$3602 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46046 \$16 \$4562 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46047 \$16 \$3691 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46051 \$153 \$4836 \$4737 \$3691 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46052 \$153 \$4738 \$4737 \$4129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46053 \$153 \$4517 \$3893 \$4857 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46055 \$153 \$4702 \$3860 \$4646 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46056 \$153 \$4647 \$4739 \$4129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46058 \$153 \$4763 \$4739 \$3826 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46059 \$16 \$4837 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46060 \$153 \$4592 \$4414 \$4371 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46061 \$16 \$3826 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46062 \$16 \$3898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46063 \$153 \$4702 \$4739 \$3898 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46064 \$16 \$3602 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46067 \$16 \$4784 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46069 \$16 \$4057 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46070 \$153 \$4290 \$3142 \$4371 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46071 \$153 \$4765 \$4739 \$4057 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46072 \$16 \$4129 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46073 \$153 \$4838 \$4740 \$4129 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46074 \$16 \$3680 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46075 \$16 \$3691 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46077 \$153 \$4764 \$4740 \$3691 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46078 \$153 \$4839 \$4740 \$3680 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46079 \$153 \$4766 \$4740 \$3602 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46080 \$16 \$3680 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46081 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$46082 \$16 \$3826 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46085 \$153 \$4840 \$4740 \$3826 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46087 \$153 \$5238 \$4740 \$3721 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46089 \$153 \$3863 \$4414 \$3899 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46090 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$46093 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$46094 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$46096 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$46097 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$46098 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$46099 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$46100 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$46101 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$46102 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$46103 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$46104 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$46107 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$46108 \$153 \$13335 \$12412 \$13336 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46109 \$153 \$13452 \$12209 \$13336 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46110 \$153 \$13399 \$12208 \$13336 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46111 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$46113 \$16 \$11757 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46114 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$46117 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$46119 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$46120 \$153 \$13453 \$12353 \$13336 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46121 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$46122 \$16 \$11757 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46123 \$153 \$13454 \$13130 \$12152 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46124 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$46127 \$153 \$13454 \$12209 \$13239 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46128 \$16 \$12152 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46129 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$46130 \$153 \$13455 \$13130 \$12230 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46131 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$46132 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$46134 \$16 \$12230 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46135 \$153 \$13455 \$12412 \$13239 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46137 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$46138 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$46139 \$153 \$13434 \$13250 \$12095 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46140 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$46141 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$46143 \$153 \$13456 \$12208 \$13369 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46145 \$153 \$13400 \$12134 \$13369 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46146 \$153 \$13484 \$13250 \$12230 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46148 \$153 \$13531 \$12134 \$13215 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46149 \$153 \$13532 \$12412 \$13215 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46152 \$153 \$13484 \$12412 \$13369 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46154 \$16 \$12230 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46155 \$16 \$13215 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46156 \$16 \$13215 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46159 \$153 \$13457 \$13115 \$12152 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46160 \$153 \$13518 \$13115 \$12236 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46161 \$16 \$12152 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46162 \$16 \$12236 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46165 \$153 \$13457 \$12209 \$13194 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46167 \$153 \$13518 \$12134 \$13194 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46169 \$153 \$13487 \$13188 \$12236 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46171 \$153 \$13519 \$13188 \$12152 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46173 \$16 \$12236 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46174 \$16 \$12152 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46175 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$46177 \$153 \$13519 \$12209 \$13216 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46178 \$153 \$13435 \$13188 \$12095 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46179 \$153 \$13487 \$12134 \$13216 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46181 \$16 \$12095 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46182 \$153 \$13458 \$12134 \$13343 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46183 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$46184 \$153 \$13488 \$13272 \$12294 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46186 \$153 \$13436 \$13272 \$12152 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46187 \$153 \$13402 \$12057 \$13343 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46188 \$153 \$13488 \$12208 \$13343 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46189 \$16 \$12294 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46192 \$153 \$13496 \$13272 \$12230 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46193 \$16 \$12152 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46196 \$153 \$13496 \$12412 \$13343 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46197 \$153 \$13532 \$13305 \$12230 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46198 \$153 \$13437 \$13305 \$12095 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46199 \$16 \$12230 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46200 \$16 \$12003 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46203 \$16 \$12230 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46205 \$16 \$12236 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46206 \$16 \$13215 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46208 \$16 \$12095 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46209 \$153 \$13533 \$13305 \$12152 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46210 \$153 \$13459 \$13305 \$12294 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46211 \$16 \$12152 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46213 \$16 \$12294 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46214 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$46215 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$46217 \$16 \$12152 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46218 \$153 \$13460 \$13298 \$12294 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46219 \$153 \$13520 \$13298 \$12152 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46220 \$153 \$13520 \$12209 \$13345 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46221 \$153 \$13460 \$12208 \$13345 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46222 \$16 \$12294 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46225 \$153 \$13497 \$13298 \$12095 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46226 \$153 \$13438 \$13298 \$12230 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46227 \$153 \$13497 \$12353 \$13345 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46228 \$16 \$12236 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46229 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$46231 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$46232 \$153 \$13489 \$12155 \$13373 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46233 \$16 \$12230 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46236 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$46238 \$153 \$13485 \$13347 \$12259 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46239 \$153 \$13489 \$13347 \$12295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46240 \$16 \$12259 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46242 \$153 \$13485 \$12307 \$13373 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46243 \$16 \$12295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46244 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$46246 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$46248 \$153 \$13498 \$13347 \$12241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46249 \$153 \$13490 \$13347 \$12160 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46252 \$153 \$13490 \$12028 \$13373 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46253 \$16 \$12160 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46254 \$16 \$12241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46255 \$16 \$13215 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46257 \$153 \$13498 \$12363 \$13373 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46258 \$16 \$12083 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46259 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$46260 \$153 \$13439 \$13220 \$12259 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46261 \$153 \$13533 \$12209 \$13215 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46263 \$16 \$12241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46265 \$153 \$13486 \$13220 \$12160 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46266 \$16 \$12259 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46267 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$46269 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$46270 \$153 \$13521 \$13220 \$12295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46271 \$153 \$13486 \$12028 \$13222 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46272 \$153 \$13521 \$12155 \$13222 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46274 \$16 \$12295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46275 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$46276 \$153 \$13499 \$13275 \$12259 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46279 \$153 \$13461 \$12028 \$13327 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46280 \$153 \$13499 \$12307 \$13327 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46281 \$16 \$12259 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46282 \$16 \$12296 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46283 \$16 \$12160 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46284 \$153 \$13491 \$13275 \$12295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46285 \$16 \$11794 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46286 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$46289 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$46291 \$153 \$13491 \$12155 \$13327 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46292 \$153 \$13389 \$13276 \$12259 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46293 \$16 \$12295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46296 \$153 \$13462 \$12363 \$13327 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46297 \$16 \$12259 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46298 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$46302 \$153 \$13464 \$13276 \$12160 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46303 \$153 \$13390 \$13276 \$12241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46304 \$153 \$13463 \$12155 \$13240 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46305 \$153 \$13464 \$12028 \$13240 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46306 \$16 \$12160 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46307 \$16 \$12241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46308 \$153 \$13500 \$13190 \$12295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46312 \$153 \$13534 \$13190 \$12241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46313 \$16 \$12295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46315 \$153 \$13500 \$12155 \$13241 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46317 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$46318 \$153 \$13440 \$13190 \$12259 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46319 \$16 \$12241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46321 \$153 \$13534 \$12363 \$13241 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46322 \$16 \$12259 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46325 \$153 \$13522 \$13224 \$12295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46326 \$153 \$13441 \$13224 \$12160 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46327 \$16 \$12295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46328 \$16 \$12160 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46330 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$46331 \$153 \$13442 \$13224 \$12241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46332 \$153 \$13492 \$13224 \$12259 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46335 \$153 \$13492 \$12307 \$13242 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46336 \$16 \$12259 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46337 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$46338 \$16 \$12241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46340 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$46342 \$153 \$13514 \$12956 \$12295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46343 \$153 \$13501 \$12956 \$12259 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46344 \$16 \$12295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46345 \$153 \$13501 \$12307 \$13051 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46346 \$153 \$13443 \$12956 \$12241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46349 \$16 \$12259 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46350 \$153 \$13523 \$13376 \$12259 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46351 \$16 \$12259 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46352 \$16 \$12160 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46353 \$16 \$12241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46354 \$16 \$11814 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46356 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$46357 \$153 \$13523 \$12307 \$13243 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46358 \$16 \$12295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46359 \$153 \$13502 \$13376 \$12295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46361 \$153 \$13465 \$12028 \$13243 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46362 \$16 \$12241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46363 \$153 \$13257 \$13376 \$12241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46364 \$153 \$13502 \$12155 \$13243 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46365 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$46366 \$153 \$13407 \$12068 \$13243 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46368 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$46369 \$16 \$12571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46370 \$153 \$13535 \$13330 \$12571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46371 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$46373 \$16 \$12297 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46375 \$153 \$13444 \$13330 \$12297 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46376 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$46378 \$16 \$12233 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46379 \$153 \$13445 \$13330 \$12233 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46380 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$46382 \$153 \$13392 \$13330 \$12298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46383 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$46384 \$16 \$12298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46385 \$16 \$12233 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46386 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$46387 \$153 \$13503 \$13258 \$12233 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46389 \$153 \$13535 \$12309 \$13244 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46391 \$153 \$13503 \$12603 \$13200 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46394 \$16 \$12297 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46395 \$153 \$13504 \$13258 \$12297 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46396 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$46398 \$16 \$12298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46399 \$153 \$13504 \$12582 \$13200 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46400 \$16 \$12571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46401 \$16 \$12233 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46402 \$153 \$13446 \$13315 \$12571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46404 \$153 \$13524 \$13315 \$12298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46405 \$153 \$13505 \$13315 \$12233 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46407 \$153 \$13524 \$12165 \$13245 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46409 \$153 \$13505 \$12603 \$13245 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46412 \$153 \$13506 \$13315 \$12297 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46413 \$153 \$13506 \$12582 \$13245 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46415 \$16 \$12297 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46417 \$16 \$12298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46418 \$153 \$13493 \$13316 \$12571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46419 \$153 \$13515 \$13316 \$12298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46421 \$153 \$13493 \$12309 \$13302 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46422 \$16 \$12233 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46423 \$153 \$13394 \$13316 \$12233 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46425 \$153 \$13355 \$12264 \$13302 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46428 \$153 \$13466 \$12582 \$13302 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46430 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$46432 \$16 \$12297 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46433 \$153 \$13467 \$13285 \$12297 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46434 \$153 \$13525 \$12165 \$13203 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46436 \$153 \$13525 \$13285 \$12298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46437 \$153 \$13467 \$12582 \$13203 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46438 \$16 \$12298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46439 \$153 \$13468 \$12309 \$13203 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46440 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$46441 \$153 \$13469 \$12603 \$13203 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46442 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$46444 \$16 \$12233 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46445 \$153 \$13526 \$13054 \$12233 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46446 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$46448 \$16 \$12297 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46450 \$153 \$13447 \$13054 \$12297 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46451 \$153 \$13526 \$12603 \$12648 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46453 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$46456 \$16 \$12571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46457 \$16 \$12298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46458 \$153 \$13507 \$13260 \$12571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46459 \$153 \$13516 \$13260 \$12298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46460 \$16 \$12297 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46461 \$153 \$13507 \$12309 \$13109 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46462 \$153 \$13448 \$13260 \$12297 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46464 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$46465 \$153 \$13431 \$12603 \$13109 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46468 \$16 \$12298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46469 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$46470 \$153 \$13536 \$13110 \$12298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46471 \$16 \$12233 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46472 \$153 \$13508 \$13110 \$12233 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46474 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$46475 \$16 \$12571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46477 \$153 \$13508 \$12603 \$13205 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46478 \$153 \$13470 \$13110 \$12571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46479 \$153 \$13536 \$12165 \$13205 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46480 \$153 \$13470 \$12309 \$13205 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46482 \$16 \$12297 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46485 \$153 \$13527 \$13395 \$12297 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46486 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$46490 \$16 \$12571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46491 \$16 \$12164 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46492 \$153 \$13411 \$12309 \$13149 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46493 \$153 \$13527 \$12582 \$13232 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46494 \$153 \$13509 \$13395 \$12164 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46497 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$46499 \$16 \$12233 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46500 \$153 \$13509 \$12217 \$13232 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46501 \$153 \$13472 \$13395 \$12233 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46502 \$153 \$13471 \$12309 \$13232 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46503 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$46504 \$153 \$13472 \$12603 \$13232 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46506 \$16 \$12287 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46507 \$153 \$13528 \$12918 \$12287 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46510 \$153 \$13449 \$12918 \$12299 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46511 \$153 \$13528 \$12339 \$13362 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46512 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$46514 \$153 \$13473 \$12918 \$12303 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46516 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$46517 \$153 \$13494 \$12918 \$12351 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46518 \$153 \$13473 \$12227 \$13362 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46519 \$16 \$12303 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46520 \$16 \$12351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46521 \$153 \$13494 \$12119 \$13362 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46522 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$46525 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$46527 \$153 \$13432 \$12119 \$13056 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46528 \$16 \$12303 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46530 \$153 \$13396 \$13094 \$12303 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46531 \$153 \$13474 \$12371 \$13056 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46532 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$46533 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$46535 \$16 \$12303 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46536 \$16 \$12351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46538 \$153 \$13495 \$13152 \$12303 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46539 \$153 \$13517 \$13152 \$12351 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46540 \$153 \$13510 \$13152 \$12287 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46541 \$153 \$13495 \$12227 \$13058 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46542 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$46544 \$153 \$13510 \$12339 \$13058 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46545 \$16 \$12287 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46548 \$16 \$12303 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46549 \$153 \$13511 \$13180 \$12303 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46550 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$46551 \$16 \$12351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46552 \$153 \$13511 \$12227 \$13181 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46553 \$16 \$12287 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46554 \$153 \$13512 \$13180 \$12287 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46556 \$153 \$13262 \$13180 \$12351 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46558 \$16 \$12303 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46559 \$153 \$13512 \$12339 \$13181 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46560 \$153 \$13476 \$13289 \$12303 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46561 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$46563 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$46566 \$153 \$13476 \$12227 \$13237 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46567 \$153 \$13477 \$12119 \$13237 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46568 \$153 \$13450 \$13289 \$12299 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46569 \$16 \$12299 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46570 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$46571 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$46573 \$153 \$13478 \$12339 \$13237 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46574 \$16 \$12287 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46575 \$153 \$13479 \$13291 \$12287 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46577 \$153 \$13433 \$13291 \$12351 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46578 \$153 \$13479 \$12339 \$13247 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46579 \$16 \$12351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46582 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$46583 \$16 \$12303 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46585 \$153 \$13480 \$13291 \$12303 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46586 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$46587 \$153 \$13480 \$12227 \$13247 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46588 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$46591 \$16 \$12287 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46592 \$153 \$13481 \$13126 \$12303 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46593 \$153 \$13529 \$13126 \$12287 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46594 \$153 \$13481 \$12227 \$13209 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46595 \$153 \$13529 \$12339 \$13209 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46596 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$46599 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$46602 \$16 \$13451 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46603 \$16 \$12010 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46604 \$16 \$13451 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46605 \$153 \$11612 \$10376 \$13451 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46606 \$16 \$13451 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46607 \$153 \$11923 \$10815 \$13451 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46608 \$153 \$13483 \$12227 \$13248 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46609 \$153 \$11791 \$10694 \$13451 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46610 \$153 \$13483 \$13156 \$12303 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46612 \$153 \$13334 \$13156 \$12287 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46613 \$16 \$12287 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46614 \$153 \$13513 \$13265 \$12287 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46615 \$16 \$12287 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46617 \$153 \$13513 \$12339 \$13249 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46619 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$46621 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$46622 \$16 \$12351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46623 \$153 \$13530 \$13265 \$12351 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46624 \$16 \$12303 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46625 \$153 \$13482 \$13265 \$12303 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46627 \$153 \$13482 \$12227 \$13249 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46628 \$16 \$13451 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46630 \$153 \$13530 \$12119 \$13249 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46631 \$153 \$11985 \$10560 \$13451 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46632 \$153 \$11852 \$10587 \$13451 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46633 \$16 \$13451 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46635 \$16 \$13451 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46636 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$46637 \$16 \$11713 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46638 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$46643 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$46644 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$46646 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$46647 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$46648 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$46649 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$46652 \$153 \$2096 \$2193 \$2006 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46653 \$153 \$2324 \$2193 \$1658 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46654 \$16 \$2006 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46655 \$16 \$1658 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46656 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$46657 \$16 \$2006 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46658 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$46660 \$153 \$2322 \$2193 \$1942 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46662 \$153 \$2111 \$2193 \$1795 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46663 \$16 \$1942 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46664 \$153 \$2351 \$1815 \$2343 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46665 \$16 \$1795 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46666 \$153 \$2274 \$2193 \$2024 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46669 \$153 \$2323 \$2193 \$2180 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46670 \$16 \$2024 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46671 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$46672 \$153 \$2415 \$2377 \$1658 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46674 \$16 \$585 \$1430 \$2352 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$46675 \$153 \$2377 \$1596 \$2352 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$46677 \$16 \$585 \$16 \$153 \$2179 VNB sky130_fd_sc_hd__inv_1
X$46678 \$153 \$2440 \$1792 \$2179 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46679 \$153 \$2378 \$1763 \$1942 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46680 \$153 \$2432 \$2210 \$2179 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46681 \$153 \$2416 \$1815 \$2179 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46682 \$16 \$1942 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46683 \$16 \$2006 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46685 \$153 \$2211 \$1763 \$2006 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46686 \$16 \$585 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46688 \$16 \$1263 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46689 \$16 \$1942 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46690 \$153 \$2441 \$1888 \$1942 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46691 \$153 \$2379 \$1888 \$2180 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46693 \$16 \$2180 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46695 \$153 \$2378 \$2064 \$1789 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46697 \$16 \$1291 \$1522 \$2353 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$46698 \$153 \$2379 \$2252 \$1861 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46699 \$153 \$2380 \$1263 \$2353 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$46700 \$153 \$2381 \$2380 \$2180 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46701 \$16 \$1522 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46702 \$16 \$1658 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46704 \$153 \$1631 \$2380 \$1658 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46705 \$16 \$1291 \$16 \$153 \$1594 VNB sky130_fd_sc_hd__inv_1
X$46706 \$16 \$2180 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46708 \$153 \$2289 \$2354 \$1980 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46709 \$16 \$1687 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46711 \$153 \$2382 \$2354 \$1687 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46713 \$153 \$2433 \$2009 \$2275 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46714 \$153 \$2383 \$2354 \$1658 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46715 \$153 \$2382 \$1792 \$2181 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46716 \$153 \$2405 \$2354 \$1795 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46717 \$16 \$1687 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46718 \$16 \$1658 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46722 \$16 \$1795 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46723 \$153 \$2139 \$2064 \$1767 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46724 \$153 \$2417 \$2252 \$2181 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46725 \$153 \$2405 \$1815 \$2181 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46726 \$153 \$2383 \$1547 \$2181 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46728 \$153 \$2325 \$2290 \$1658 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46729 \$16 \$2442 \$16 \$153 \$1430 VNB sky130_fd_sc_hd__clkbuf_2
X$46731 \$153 \$2443 \$2290 \$2180 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46732 \$153 \$2325 \$1547 \$2344 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46734 \$16 \$849 \$16 \$153 \$2344 VNB sky130_fd_sc_hd__inv_1
X$46735 \$153 \$2381 \$2252 \$1594 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46736 \$153 \$2418 \$2290 \$1942 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46738 \$153 \$2384 \$2290 \$1687 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46740 \$153 \$2384 \$1792 \$2344 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46742 \$153 \$2291 \$2194 \$2024 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46743 \$153 \$2418 \$2064 \$2344 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46746 \$16 \$849 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46747 \$16 \$1594 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46748 \$153 \$2385 \$2194 \$1942 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46750 \$153 \$2444 \$2478 \$1942 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46751 \$16 \$2024 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46752 \$16 \$1942 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46753 \$16 \$2180 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46754 \$16 \$1942 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46755 \$16 \$2006 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46757 \$16 \$2180 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46761 \$153 \$2217 \$1792 \$2219 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46762 \$153 \$2292 \$2252 \$2219 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46763 \$153 \$2477 \$2252 \$2386 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46764 \$16 \$1596 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46765 \$153 \$2293 \$1943 \$2219 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46766 \$153 \$2444 \$2064 \$2386 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46767 \$16 \$716 \$16 \$153 \$2386 VNB sky130_fd_sc_hd__inv_1
X$46768 \$153 \$2326 \$2194 \$1980 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46771 \$153 \$2478 \$584 \$2419 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$46772 \$153 \$2326 \$2009 \$2219 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46773 \$16 \$716 \$2647 \$2419 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$46776 \$16 \$2445 \$16 \$153 \$1037 VNB sky130_fd_sc_hd__clkbuf_2
X$46777 \$16 \$2387 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46778 \$16 \$2387 \$16 \$153 \$2183 VNB sky130_fd_sc_hd__clkbuf_2
X$46779 \$153 \$2182 \$2420 \$2435 \$2436 \$2434 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4bb_2
X$46781 \$16 \$2220 \$2196 \$2183 \$153 \$2114 \$16 VNB sky130_fd_sc_hd__and3b_4
X$46782 \$16 \$2233 \$16 \$153 \$2220 VNB sky130_fd_sc_hd__clkbuf_2
X$46783 \$16 \$2183 \$2220 \$2196 \$153 \$16 \$2276 VNB sky130_fd_sc_hd__and3_4
X$46784 \$16 \$2233 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46785 \$153 \$2296 \$2434 \$2436 \$2420 \$2435 \$16 \$16 VNB
+ sky130_fd_sc_hd__nor4b_2
X$46786 \$16 \$1354 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46788 \$153 \$2389 \$1596 \$2295 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$46789 \$16 \$2675 \$16 \$153 \$1480 VNB sky130_fd_sc_hd__clkbuf_2
X$46791 \$16 \$1923 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46792 \$153 \$2388 \$1895 \$2390 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46793 \$153 \$2388 \$2389 \$1923 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46794 \$153 \$2421 \$2184 \$2390 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46795 \$153 \$2481 \$1806 \$2390 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46796 \$16 \$2355 \$16 \$153 \$716 VNB sky130_fd_sc_hd__clkbuf_2
X$46798 \$16 \$2356 \$16 \$153 \$1551 VNB sky130_fd_sc_hd__clkbuf_2
X$46800 \$153 \$2446 \$2389 \$2042 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46801 \$16 \$2199 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46802 \$153 \$2297 \$2026 \$1944 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46803 \$16 \$585 \$16 \$153 \$2390 VNB sky130_fd_sc_hd__inv_1
X$46804 \$153 \$2447 \$2026 \$2390 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46806 \$153 \$2116 \$2039 \$1805 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46809 \$153 \$2437 \$2389 \$1845 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46810 \$153 \$2357 \$1954 \$2390 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46811 \$153 \$2391 \$1703 \$2390 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46812 \$16 \$1845 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46813 \$16 \$2634 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46814 \$153 \$2406 \$2244 \$2042 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46815 \$16 \$2634 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46818 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$46820 \$16 \$1805 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46821 \$153 \$2392 \$2244 \$1965 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46822 \$153 \$2437 \$1471 \$2390 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46823 \$153 \$2448 \$2026 \$2299 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46824 \$153 \$2393 \$2244 \$1923 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46825 \$16 \$2042 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46827 \$153 \$2392 \$1806 \$2299 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46829 \$153 \$2449 \$1921 \$2199 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46830 \$153 \$2394 \$1921 \$2042 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46831 \$153 \$2394 \$1924 \$1922 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46834 \$16 \$2042 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46835 \$16 \$1291 \$1966 \$2358 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$46836 \$153 \$2359 \$1263 \$2358 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$46837 \$153 \$2300 \$1471 \$1922 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46838 \$16 \$2199 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46840 \$153 \$2450 \$1471 \$2327 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46841 \$16 \$1263 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46842 \$16 \$1291 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46843 \$153 \$2301 \$2184 \$1866 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46845 \$153 \$2360 \$2359 \$1965 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46846 \$16 \$1291 \$16 \$153 \$2327 VNB sky130_fd_sc_hd__inv_1
X$46847 \$153 \$2360 \$1806 \$2327 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46848 \$16 \$1965 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46849 \$153 \$2361 \$1924 \$2327 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46851 \$153 \$2277 \$1047 \$2223 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$46854 \$16 \$2362 \$16 \$153 \$1966 VNB sky130_fd_sc_hd__clkbuf_2
X$46855 \$16 \$1966 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46856 \$16 \$1067 \$1966 \$2451 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$46857 \$16 \$1067 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46858 \$153 \$2328 \$2277 \$2043 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46860 \$153 \$2345 \$2277 \$2199 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46861 \$16 \$2043 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46862 \$153 \$2328 \$1954 \$2152 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46865 \$153 \$2452 \$2184 \$2499 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46866 \$153 \$2345 \$2184 \$2152 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46867 \$16 \$2199 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46868 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$46869 \$153 \$2422 \$2277 \$1923 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46871 \$16 \$1659 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46872 \$153 \$2363 \$1471 \$2346 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46875 \$16 \$1965 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46876 \$153 \$2422 \$1895 \$2152 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46877 \$153 \$2200 \$1659 \$2329 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$46878 \$16 \$1923 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46879 \$16 \$1966 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46880 \$16 \$899 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46881 \$16 \$1845 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46882 \$153 \$2330 \$2200 \$1965 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46883 \$153 \$2225 \$1895 \$2186 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46885 \$16 \$899 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46887 \$153 \$2453 \$2184 \$2186 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46889 \$153 \$2395 \$2200 \$2042 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46890 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$46891 \$16 \$716 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46892 \$16 \$2042 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46893 \$153 \$2395 \$1924 \$2186 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46895 \$16 \$716 \$2347 \$2396 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$46898 \$153 \$2454 \$1703 \$2186 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46899 \$153 \$2365 \$584 \$2396 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$46900 \$16 \$652 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46901 \$153 \$2119 \$2365 \$1923 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46902 \$16 \$652 \$2347 \$2302 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$46904 \$153 \$2397 \$2365 \$1805 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46906 \$16 \$716 \$16 \$153 \$2120 VNB sky130_fd_sc_hd__inv_1
X$46907 \$16 \$1923 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46909 \$153 \$2397 \$1703 \$2120 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46910 \$16 \$1805 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46912 \$153 \$2331 \$2365 \$2089 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46914 \$153 \$2408 \$2365 \$1965 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46916 \$16 \$2089 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46917 \$16 \$1845 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46918 \$153 \$2455 \$2365 \$1845 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46919 \$153 \$2331 \$2026 \$2120 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46920 \$153 \$2408 \$1806 \$2120 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46921 \$16 \$1965 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46922 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$46924 \$153 \$2366 \$2279 \$2098 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46926 \$153 \$2456 \$2279 \$1879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46927 \$153 \$2076 \$1715 \$1540 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46928 \$16 \$1879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46930 \$16 \$594 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46931 \$16 \$2098 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46932 \$16 \$1969 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46933 \$16 \$2105 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46934 \$153 \$2423 \$2279 \$2105 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46935 \$16 \$558 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46936 \$16 \$1878 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46938 \$153 \$2366 \$1993 \$2278 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46939 \$16 \$594 \$1968 \$2304 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$46940 \$16 \$2104 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46941 \$153 \$2423 \$2438 \$2278 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46942 \$153 \$2332 \$2279 \$2104 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46943 \$16 \$2104 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46944 \$16 \$594 \$16 \$153 \$2278 VNB sky130_fd_sc_hd__inv_1
X$46947 \$153 \$2398 \$1715 \$2278 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46948 \$153 \$2398 \$2279 \$2016 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46949 \$153 \$2409 \$2103 \$2104 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46951 \$153 \$2305 \$1715 \$2078 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46952 \$153 \$2260 \$1993 \$2078 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46954 \$153 \$2409 \$2092 \$2078 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46956 \$16 \$1756 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46957 \$153 \$2306 \$2103 \$1756 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46958 \$16 \$594 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46959 \$153 \$2077 \$1715 \$1679 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46961 \$16 \$438 \$1968 \$2457 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$46962 \$153 \$2348 \$2103 \$1969 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46963 \$16 \$438 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46965 \$16 \$438 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46966 \$16 \$884 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46967 \$16 \$964 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46968 \$16 \$2016 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46969 \$153 \$2424 \$2202 \$2016 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46970 \$153 \$2348 \$1613 \$2078 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46971 \$16 \$964 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46972 \$16 \$354 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46973 \$16 \$1628 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46974 \$16 \$1879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46975 \$153 \$2424 \$1715 \$2280 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46977 \$153 \$2307 \$1712 \$2280 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$46979 \$16 \$1878 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46980 \$153 \$2308 \$2202 \$1879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46981 \$153 \$2458 \$2202 \$1878 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46982 \$16 \$354 \$16 \$153 \$2280 VNB sky130_fd_sc_hd__inv_1
X$46983 \$16 \$1879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46984 \$16 \$674 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46986 \$16 \$2105 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46987 \$16 \$1878 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46989 \$153 \$2333 \$2309 \$1878 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46990 \$153 \$2459 \$2309 \$1879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46991 \$16 \$1811 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46992 \$16 \$1811 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46994 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$46995 \$16 \$1756 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$46996 \$153 \$2367 \$2309 \$1756 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$46998 \$153 \$2333 \$1868 \$2334 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47000 \$153 \$2367 \$1712 \$2334 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47001 \$153 \$2460 \$1715 \$2334 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47002 \$16 \$829 \$16 \$153 \$2334 VNB sky130_fd_sc_hd__inv_1
X$47003 \$16 \$1756 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47004 \$153 \$2230 \$2310 \$1756 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47005 \$16 \$829 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47006 \$16 \$2098 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47008 \$153 \$2410 \$2310 \$2098 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47010 \$153 \$2410 \$1993 \$2187 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47012 \$16 \$80 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47014 \$16 \$2104 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47015 \$16 \$1929 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47016 \$16 \$80 \$1929 \$2311 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$47017 \$153 \$2425 \$2310 \$2104 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47019 \$153 \$2263 \$1868 \$2187 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47020 \$153 \$2399 \$1715 \$2187 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47021 \$153 \$2461 \$2310 \$1879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47022 \$153 \$2312 \$1613 \$2187 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47023 \$16 \$2105 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47024 \$16 \$80 \$16 \$153 \$2187 VNB sky130_fd_sc_hd__inv_1
X$47026 \$153 \$2426 \$2368 \$2105 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47027 \$153 \$2335 \$2368 \$2016 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47028 \$153 \$2426 \$2438 \$2188 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47029 \$153 \$2335 \$1715 \$2188 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47031 \$16 \$2098 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47035 \$153 \$2336 \$2368 \$2098 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47036 \$16 \$1811 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47037 \$16 \$1878 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47038 \$153 \$2281 \$2368 \$1878 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47039 \$153 \$2336 \$1993 \$2188 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47040 \$16 \$508 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47041 \$16 \$508 \$16 \$153 \$2188 VNB sky130_fd_sc_hd__inv_1
X$47042 \$16 \$724 \$2580 \$2313 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$47043 \$16 \$2580 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47045 \$16 \$2580 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47046 \$153 \$2732 \$1600 \$2369 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$47048 \$16 \$276 \$2580 \$2369 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$47049 \$16 \$2580 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47050 \$16 \$276 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47052 \$16 \$1378 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47053 \$16 \$1600 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47054 \$16 \$2387 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47055 \$16 \$2349 \$2370 \$2315 \$153 \$2055 \$16 VNB sky130_fd_sc_hd__and3b_4
X$47056 \$16 \$1378 \$16 \$153 \$2370 VNB sky130_fd_sc_hd__clkbuf_2
X$47057 \$16 \$2387 \$16 \$153 \$2349 VNB sky130_fd_sc_hd__clkbuf_2
X$47058 \$16 \$2315 \$2370 \$2349 \$153 \$2463 \$16 VNB sky130_fd_sc_hd__and3b_4
X$47060 \$153 \$2315 \$2349 \$2400 \$2370 \$16 \$16 VNB sky130_fd_sc_hd__nor3b_4
X$47061 \$16 \$2126 \$16 \$153 \$2372 VNB sky130_fd_sc_hd__clkbuf_2
X$47062 \$16 \$2400 \$16 \$153 \$2464 VNB sky130_fd_sc_hd__clkbuf_2
X$47065 \$153 \$2439 \$2371 \$2372 \$2337 \$2464 \$16 \$16 VNB
+ sky130_fd_sc_hd__nor4b_2
X$47066 \$16 \$594 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47067 \$153 \$2372 \$2337 \$2350 \$2371 \$2464 \$16 \$16 VNB
+ sky130_fd_sc_hd__and4b_2
X$47068 \$16 \$2350 \$16 \$153 \$724 VNB sky130_fd_sc_hd__clkbuf_2
X$47070 \$16 \$2439 \$16 \$153 \$1228 VNB sky130_fd_sc_hd__clkbuf_2
X$47071 \$16 \$558 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47072 \$16 \$2465 \$16 \$153 \$276 VNB sky130_fd_sc_hd__clkbuf_2
X$47074 \$16 \$1972 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47075 \$153 \$2401 \$2316 \$2191 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47076 \$16 \$902 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47078 \$153 \$2466 \$2316 \$2031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47079 \$16 \$594 \$16 \$153 \$2402 VNB sky130_fd_sc_hd__inv_1
X$47082 \$153 \$2338 \$2316 \$2093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47083 \$153 \$2401 \$2267 \$2402 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47085 \$153 \$2374 \$2316 \$2192 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47086 \$153 \$2373 \$2316 \$1960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47087 \$16 \$2192 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47089 \$16 \$399 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47090 \$16 \$1960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47091 \$153 \$2373 \$2086 \$2402 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47092 \$16 \$2191 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47093 \$153 \$2427 \$1935 \$2191 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47094 \$153 \$2374 \$2269 \$2402 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47095 \$16 \$399 \$16 \$153 \$2506 VNB sky130_fd_sc_hd__inv_1
X$47096 \$153 \$2427 \$2267 \$2506 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47097 \$16 \$265 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47100 \$153 \$2317 \$2271 \$2129 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47102 \$153 \$2411 \$1935 \$2093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47104 \$153 \$2170 \$1936 \$2129 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47105 \$153 \$2411 \$2265 \$2506 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47106 \$16 \$438 \$1972 \$2467 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$47107 \$16 \$1972 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47110 \$16 \$2191 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47111 \$16 \$438 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47112 \$153 \$2339 \$1909 \$2191 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47114 \$153 \$2428 \$1909 \$2192 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47116 \$153 \$2339 \$2267 \$1870 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47117 \$153 \$2428 \$2269 \$1870 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47119 \$16 \$2192 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47120 \$153 \$2318 \$2271 \$1870 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47121 \$16 \$2031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47122 \$16 \$1960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47123 \$153 \$2340 \$2099 \$1960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47125 \$16 \$2085 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47126 \$153 \$2429 \$2099 \$2085 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47127 \$153 \$2340 \$2086 \$2239 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47130 \$153 \$2429 \$2271 \$2239 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47131 \$16 \$2192 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47132 \$153 \$2341 \$2099 \$2192 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47134 \$16 \$2191 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47135 \$153 \$2412 \$2099 \$2191 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47137 \$16 \$80 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47138 \$16 \$116 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47139 \$16 \$2093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47142 \$153 \$2412 \$2267 \$2239 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47143 \$153 \$2468 \$2099 \$2093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47144 \$153 \$2403 \$116 \$2375 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$47145 \$16 \$80 \$1885 \$2375 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$47147 \$16 \$724 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47148 \$16 \$1885 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47149 \$16 \$2085 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47150 \$16 \$1860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47151 \$153 \$2319 \$1886 \$2085 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47153 \$153 \$2469 \$2403 \$1860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47154 \$153 \$2493 \$2056 \$2282 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47155 \$16 \$80 \$16 \$153 \$2282 VNB sky130_fd_sc_hd__inv_1
X$47157 \$153 \$2413 \$2403 \$2031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47159 \$16 \$1960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47161 \$153 \$2283 \$2403 \$1960 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47163 \$16 \$276 \$2531 \$2430 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$47164 \$153 \$2376 \$1600 \$2430 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$47165 \$153 \$2413 \$1936 \$2282 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47166 \$16 \$2085 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47167 \$16 \$2093 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47169 \$153 \$2342 \$2376 \$2093 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47170 \$153 \$2320 \$2376 \$2085 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47172 \$153 \$2342 \$2265 \$2284 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47173 \$153 \$2431 \$2376 \$2191 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47174 \$16 \$2191 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47176 \$153 \$2404 \$2376 \$1860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47177 \$153 \$2431 \$2267 \$2284 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47178 \$153 \$2404 \$2000 \$2284 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47179 \$153 \$2285 \$2376 \$1973 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47180 \$16 \$1973 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47182 \$16 \$2031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47185 \$16 \$1960 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47188 \$153 \$2321 \$2376 \$2192 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47189 \$153 \$2208 \$2376 \$2031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47190 \$153 \$2273 \$2086 \$2284 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47191 \$16 \$2192 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47192 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$47195 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$47196 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$47198 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$47199 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$47200 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$47201 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$47202 \$153 \$6708 \$3284 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$47203 \$16 \$6708 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47204 \$16 \$6783 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47205 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$47206 \$153 \$6730 \$6403 \$5518 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47207 \$16 \$5518 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47208 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$47210 \$153 \$6603 \$5373 \$6452 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47211 \$153 \$6730 \$5463 \$6452 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47213 \$153 \$6661 \$5373 \$6257 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47214 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$47215 \$153 \$6662 \$5463 \$6257 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47216 \$153 \$6717 \$6719 \$6709 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47219 \$153 \$6691 \$6251 \$5489 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47220 \$153 \$6731 \$6782 \$6860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47221 \$16 \$5489 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47222 \$16 \$6860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47224 \$153 \$6604 \$5177 \$6315 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47225 \$153 \$6663 \$5373 \$6315 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47229 \$153 \$6664 \$5174 \$6315 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47230 \$153 \$6718 \$6719 \$6815 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47231 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$47232 \$153 \$6665 \$5373 \$6409 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47233 \$153 \$6720 \$6732 \$6815 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47234 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$47235 \$153 \$6819 \$6719 \$6692 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47238 \$16 \$6733 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47239 \$16 \$6900 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47241 \$16 \$6693 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47242 \$153 \$6721 \$6732 \$6692 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47243 \$153 \$6693 \$3333 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$47244 \$153 \$6666 \$3491 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$47246 \$153 \$6694 \$6341 \$5489 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47247 \$153 \$6694 \$5373 \$6316 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47249 \$153 \$6820 \$3335 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$47250 \$153 \$6607 \$5463 \$6316 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47253 \$153 \$6722 \$3244 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$47254 \$153 \$6766 \$6749 \$6857 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47255 \$153 \$6822 \$6749 \$6710 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47256 \$153 \$6723 \$7003 \$6711 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47257 \$153 \$6724 \$6732 \$6710 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47259 \$153 \$6712 \$3096 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$47260 \$16 \$5518 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47261 \$16 \$3096 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47262 \$153 \$6570 \$6435 \$5467 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47263 \$16 \$5467 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47264 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$47266 \$153 \$6668 \$5390 \$6453 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47268 \$153 \$6734 \$6435 \$5566 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47270 \$153 \$6799 \$1918 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$47271 \$153 \$6541 \$5287 \$6453 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47272 \$153 \$6725 \$6906 \$6695 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47275 \$153 \$6726 \$6906 \$6713 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47276 \$153 \$6669 \$1775 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$47277 \$16 \$5478 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47278 \$153 \$6576 \$6326 \$5478 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47279 \$153 \$6463 \$5406 \$6264 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47281 \$153 \$6625 \$5205 \$6264 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47282 \$16 \$5478 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47284 \$153 \$6577 \$6440 \$5566 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47285 \$153 \$6696 \$6440 \$5478 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47286 \$153 \$6696 \$5390 \$6357 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47287 \$16 \$5478 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47289 \$153 \$6578 \$6344 \$5478 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47290 \$16 \$5478 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47292 \$16 \$6797 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47294 \$153 \$6579 \$6344 \$5566 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47295 \$153 \$6670 \$5205 \$6358 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47296 \$16 \$5566 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47297 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$47299 \$16 \$6735 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47301 \$153 \$6735 \$1406 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$47302 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$47303 \$153 \$6580 \$6034 \$5478 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47304 \$153 \$6672 \$5205 \$6291 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47305 \$16 \$5478 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47308 \$153 \$6611 \$5406 \$6291 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47309 \$16 \$6754 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47311 \$153 \$3508 \$5478 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$47313 \$153 \$3243 \$5232 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$47315 \$16 \$1406 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47317 \$153 \$1406 \$5605 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$47319 \$16 \$5932 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47320 \$16 \$5819 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47321 \$16 \$1918 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47322 \$153 \$1918 \$5834 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$47323 \$153 \$6727 \$6200 \$6556 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47325 \$153 \$6697 \$6642 \$5528 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47327 \$153 \$6736 \$6698 \$5528 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47328 \$16 \$5528 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47330 \$153 \$6698 \$5480 \$6615 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$47331 \$16 \$5480 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47332 \$16 \$5702 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47333 \$16 \$4834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47335 \$153 \$6673 \$6200 \$6616 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47336 \$16 \$5819 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47337 \$153 \$6737 \$6585 \$5819 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47339 \$153 \$6699 \$6585 \$5796 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47340 \$153 \$6699 \$5775 \$6617 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47341 \$16 \$5819 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47345 \$16 \$5834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47346 \$153 \$6674 \$6200 \$6714 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47347 \$153 \$6700 \$6643 \$5834 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47348 \$153 \$6700 \$5881 \$6714 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47350 \$16 \$5796 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47351 \$153 \$6701 \$6511 \$5796 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47353 \$153 \$6701 \$5775 \$6558 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47354 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$47355 \$16 \$5796 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47356 \$153 \$6738 \$6563 \$5796 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47357 \$16 \$5528 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47358 \$153 \$6739 \$6563 \$5528 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47359 \$16 \$5605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47360 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$47361 \$16 \$5819 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47363 \$153 \$6740 \$6645 \$5819 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47364 \$153 \$6741 \$6645 \$5528 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47365 \$16 \$5528 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47366 \$16 \$5528 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47367 \$16 \$5856 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47368 \$153 \$6702 \$6742 \$5528 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47369 \$16 \$5834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47371 \$153 \$6702 \$5500 \$6715 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47372 \$153 \$6878 \$5755 \$6715 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47374 \$153 \$6703 \$5306 \$6676 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$47375 \$153 \$6742 \$5235 \$6759 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$47376 \$153 \$6843 \$5881 \$6677 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47378 \$153 \$6743 \$6703 \$5528 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47379 \$16 \$1488 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47380 \$153 \$1488 \$5579 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$47381 \$16 \$5718 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47382 \$153 \$6704 \$6679 \$5887 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47384 \$16 \$5887 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47385 \$153 \$6704 \$5627 \$6657 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47386 \$153 \$6744 \$6679 \$5579 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47387 \$16 \$5786 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47388 \$16 \$5541 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47390 \$16 \$5579 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47391 \$153 \$6658 \$6681 \$5579 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47392 \$16 \$5351 \$16 \$153 \$6682 VNB sky130_fd_sc_hd__inv_1
X$47393 \$16 \$5351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47396 \$16 \$5786 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47397 \$153 \$6705 \$6681 \$5786 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47398 \$153 \$6705 \$5635 \$6682 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47400 \$153 \$6716 \$6619 \$5579 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47401 \$153 \$6716 \$5484 \$6639 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47402 \$16 \$5379 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47404 \$16 \$5331 \$6216 \$6683 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$47405 \$153 \$6745 \$6631 \$5579 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47406 \$153 \$6706 \$6631 \$5718 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47407 \$153 \$6706 \$5938 \$6633 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47409 \$153 \$5336 \$3986 \$4954 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47411 \$153 \$6746 \$6640 \$5718 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47412 \$153 \$6746 \$5938 \$6684 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47413 \$153 \$6564 \$6620 \$5718 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47414 \$16 \$5579 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47415 \$153 \$6685 \$5627 \$6565 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47416 \$16 \$5718 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47417 \$16 \$4803 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47419 \$16 \$5718 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47420 \$153 \$6599 \$6686 \$5718 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47422 \$153 \$6687 \$5484 \$6561 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47424 \$153 \$6707 \$6688 \$5718 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47425 \$153 \$6707 \$5938 \$6601 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47426 \$16 \$5579 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47428 \$153 \$6747 \$5235 \$6728 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$47429 \$153 \$6729 \$5484 \$6601 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47430 \$153 \$6689 \$5484 \$6457 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47431 \$16 \$5235 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47432 \$16 \$5609 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47433 \$153 \$6748 \$6562 \$5609 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47434 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$47436 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$47437 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$47438 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$47439 \$153 \$6761 \$6859 \$6783 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47441 \$153 \$6539 \$5055 \$6452 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47443 \$153 \$6477 \$5107 \$6452 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47444 \$16 \$6784 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47445 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$47446 \$153 \$6811 \$6859 \$6792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47448 \$153 \$6812 \$6781 \$6784 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47449 \$16 \$6784 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47450 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$47452 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$47453 \$153 \$6762 \$6781 \$6783 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47454 \$153 \$6762 \$6749 \$6709 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47456 \$153 \$6750 \$6782 \$6784 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47457 \$153 \$6763 \$6732 \$6709 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47460 \$153 \$6814 \$6782 \$6783 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47461 \$16 \$6783 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47462 \$153 \$6816 \$6751 \$6783 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47463 \$16 \$6783 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47464 \$153 \$6817 \$6751 \$6784 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47465 \$16 \$6784 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47468 \$153 \$6818 \$6752 \$6784 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47470 \$16 \$6792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47471 \$16 \$6784 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47472 \$16 \$6907 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47473 \$153 \$6764 \$6752 \$6783 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47474 \$153 \$6764 \$6749 \$6692 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47475 \$16 \$6783 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47476 \$16 \$6860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47477 \$16 \$6761 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47478 \$16 \$6733 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47480 \$153 \$6793 \$6794 \$6914 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47481 \$153 \$6933 \$6719 \$6914 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47482 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$47484 \$16 \$5489 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47485 \$153 \$6765 \$6785 \$6784 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47486 \$153 \$6765 \$6794 \$6795 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47487 \$16 \$6783 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47488 \$16 \$6820 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47489 \$16 \$6784 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47491 \$16 \$6753 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47492 \$16 \$7535 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47493 \$16 \$7535 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47495 \$153 \$6821 \$6786 \$6784 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47496 \$16 \$6784 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47497 \$16 \$6722 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47499 \$16 \$6783 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47500 \$153 \$6766 \$6786 \$6783 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47501 \$16 \$7041 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47502 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$47504 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$47506 \$153 \$6823 \$6861 \$6784 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47507 \$16 \$6784 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47509 \$153 \$6609 \$5463 \$6177 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47510 \$153 \$6824 \$6796 \$6797 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47511 \$16 \$6797 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47514 \$153 \$6798 \$6756 \$6711 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47515 \$153 \$6825 \$6796 \$6771 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47516 \$153 \$6734 \$5519 \$6453 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47517 \$153 \$6767 \$6787 \$6754 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47518 \$16 \$6799 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47519 \$16 \$5566 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47520 \$16 \$6754 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47522 \$16 \$6797 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47523 \$16 \$6771 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47524 \$16 \$6695 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47525 \$16 \$6695 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47526 \$153 \$6726 \$6755 \$6797 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47527 \$16 \$5566 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47529 \$153 \$6768 \$6755 \$6754 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47530 \$153 \$6768 \$6756 \$6713 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47531 \$16 \$6754 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47532 \$16 \$6695 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47534 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$47535 \$153 \$6800 \$6865 \$6652 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47536 \$153 \$6769 \$6326 \$5566 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47537 \$153 \$6769 \$5519 \$6264 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47538 \$16 \$5566 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47540 \$153 \$6770 \$6788 \$6771 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47542 \$153 \$6770 \$6865 \$6801 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47543 \$16 \$5566 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47544 \$16 \$6771 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47545 \$16 \$6754 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47546 \$153 \$6827 \$6788 \$6754 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47547 \$153 \$6828 \$6788 \$6797 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47548 \$153 \$6829 \$6867 \$6803 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47551 \$153 \$6830 \$6789 \$6797 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47552 \$153 \$6802 \$6865 \$6803 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47553 \$16 \$6797 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47555 \$153 \$6772 \$6790 \$6754 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47556 \$153 \$6804 \$7003 \$6805 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47557 \$16 \$6754 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47559 \$153 \$6831 \$6790 \$6771 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47561 \$153 \$6893 \$1407 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$47562 \$153 \$6773 \$6791 \$6754 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47564 \$16 \$6771 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47566 \$153 \$6832 \$6791 \$6771 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47567 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$47569 \$16 \$1407 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47570 \$153 \$1407 \$5714 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$47572 \$16 \$5819 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47573 \$153 \$6806 \$5775 \$6556 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47575 \$153 \$6727 \$6642 \$5819 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47576 \$153 \$6655 \$6642 \$5834 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47577 \$16 \$5714 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47578 \$16 \$5528 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47579 \$16 \$5856 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47580 \$16 \$5856 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47581 \$153 \$6636 \$6698 \$5714 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47583 \$16 \$5351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47584 \$153 \$6736 \$5500 \$6616 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47585 \$16 \$5834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47586 \$153 \$6757 \$6698 \$5834 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47588 \$16 \$5834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47589 \$153 \$6834 \$6585 \$5834 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47590 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$47592 \$16 \$5796 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47594 \$153 \$6737 \$6200 \$6617 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47595 \$153 \$6947 \$5470 \$6617 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47597 \$16 \$5714 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47598 \$153 \$6758 \$6643 \$5714 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47599 \$153 \$6675 \$5500 \$6714 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47600 \$153 \$6758 \$5755 \$6714 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47603 \$16 \$5331 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47604 \$16 \$5331 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47605 \$16 \$5834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47606 \$153 \$6774 \$6511 \$5834 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47607 \$16 \$6656 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47608 \$153 \$6774 \$5881 \$6558 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47609 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$47610 \$16 \$5714 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47611 \$16 \$5856 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47612 \$153 \$6775 \$6563 \$5714 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47614 \$153 \$6738 \$5775 \$6533 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47616 \$153 \$6739 \$5500 \$6533 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47617 \$153 \$6839 \$6645 \$5605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47618 \$153 \$6740 \$6200 \$6560 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47619 \$153 \$6840 \$5775 \$6560 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47620 \$16 \$4803 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47622 \$153 \$6776 \$5881 \$6560 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47623 \$153 \$6741 \$5500 \$6560 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47624 \$153 \$6841 \$6742 \$5834 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47625 \$153 \$6842 \$6742 \$5819 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47626 \$16 \$5173 \$6269 \$6759 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$47629 \$153 \$6844 \$6703 \$5819 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47630 \$16 \$5819 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47631 \$16 \$5714 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47632 \$16 \$5528 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47633 \$153 \$6777 \$6703 \$5714 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47634 \$153 \$6743 \$5500 \$6677 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47635 \$153 \$6777 \$5755 \$6677 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47637 \$153 \$6678 \$5775 \$6535 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47639 \$16 \$5767 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47640 \$153 \$6778 \$6679 \$5767 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47641 \$153 \$6778 \$5575 \$6657 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47642 \$16 \$5579 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47643 \$153 \$6846 \$6679 \$5786 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47646 \$153 \$6744 \$5484 \$6657 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47648 \$16 \$5887 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47649 \$153 \$6847 \$6681 \$5887 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47650 \$16 \$5718 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47651 \$153 \$6659 \$6681 \$5718 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47652 \$153 \$6847 \$5627 \$6682 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47656 \$153 \$6660 \$6619 \$5718 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47657 \$153 \$6807 \$5627 \$6639 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47658 \$16 \$5718 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47660 \$16 \$5887 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47661 \$16 \$5579 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47663 \$153 \$6850 \$6631 \$5887 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47664 \$16 \$5718 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47665 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$47667 \$153 \$6745 \$5484 \$6633 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47668 \$16 \$5887 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47669 \$16 \$5579 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47670 \$153 \$6402 \$5938 \$6924 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47671 \$153 \$6808 \$6640 \$5579 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47672 \$153 \$6808 \$5484 \$6684 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47673 \$153 \$6852 \$5627 \$6684 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47675 \$153 \$6779 \$6620 \$5579 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47676 \$153 \$6779 \$5484 \$6565 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47678 \$16 \$5609 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47679 \$153 \$6780 \$6686 \$5609 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47680 \$153 \$6780 \$5074 \$6561 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47681 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$47683 \$16 \$5718 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47685 \$153 \$6809 \$5484 \$6760 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47686 \$153 \$6810 \$5627 \$6601 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47687 \$153 \$6729 \$6688 \$5579 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47688 \$153 \$6809 \$6747 \$5579 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47689 \$16 \$5173 \$16 \$153 \$6760 VNB sky130_fd_sc_hd__inv_1
X$47691 \$153 \$6554 \$5575 \$6457 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47692 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$47693 \$153 \$6372 \$5074 \$6274 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47694 \$153 \$6496 \$5627 \$6274 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47695 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$47696 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$47697 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$47698 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$47699 \$16 \$7041 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47700 \$153 \$6856 \$6930 \$6855 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47701 \$153 \$6883 \$6859 \$6784 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47702 \$153 \$6863 \$6859 \$6860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47703 \$16 \$6860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47704 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$47706 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$47707 \$16 \$6792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47709 \$153 \$6717 \$6781 \$6792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47710 \$153 \$6812 \$6794 \$6709 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47711 \$16 \$6792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47712 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$47713 \$153 \$6763 \$6781 \$6860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47714 \$16 \$6783 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47715 \$16 \$6860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47718 \$16 \$6813 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47719 \$153 \$6864 \$6782 \$6792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47720 \$153 \$6750 \$6794 \$6980 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47721 \$16 \$6792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47723 \$153 \$6814 \$6749 \$6980 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47724 \$153 \$6720 \$6751 \$6860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47726 \$16 \$6860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47727 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$47728 \$153 \$6816 \$6749 \$6815 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47729 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$47730 \$153 \$6817 \$6794 \$6815 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47731 \$153 \$6819 \$6752 \$6792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47732 \$153 \$6818 \$6794 \$6692 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47735 \$153 \$6721 \$6752 \$6860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47736 \$153 \$6793 \$6908 \$6784 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47737 \$16 \$6784 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47739 \$153 \$6884 \$6908 \$6783 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47740 \$16 \$6783 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47741 \$16 \$6860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47744 \$153 \$6885 \$6785 \$6783 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47745 \$153 \$6648 \$6785 \$6860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47746 \$16 \$6860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47747 \$16 \$6935 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47748 \$153 \$6886 \$6786 \$6860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47749 \$16 \$6860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47750 \$16 \$6887 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47752 \$153 \$6821 \$6794 \$6857 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47754 \$16 \$6783 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47755 \$153 \$6822 \$6861 \$6783 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47756 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$47757 \$153 \$6724 \$6861 \$6860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47758 \$16 \$6860 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47759 \$16 \$6888 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47760 \$16 \$6988 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47764 \$153 \$6723 \$6796 \$6862 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47765 \$153 \$6798 \$6796 \$6754 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47766 \$16 \$6754 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47767 \$153 \$6866 \$6796 \$6916 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47768 \$16 \$6916 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47769 \$16 \$6771 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47771 \$16 \$7044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47772 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$47773 \$153 \$6725 \$6787 \$6797 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47774 \$153 \$6825 \$6865 \$6711 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47775 \$153 \$6866 \$6867 \$6711 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47776 \$153 \$6767 \$6756 \$6695 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47777 \$16 \$6862 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47778 \$16 \$6797 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47781 \$153 \$6889 \$6755 \$6862 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47782 \$153 \$6868 \$6865 \$6713 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47783 \$16 \$6862 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47785 \$153 \$6826 \$6869 \$6754 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47786 \$16 \$6754 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47787 \$153 \$6826 \$6756 \$6652 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47789 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$47790 \$153 \$6890 \$6870 \$6797 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47791 \$153 \$6871 \$6865 \$6918 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47792 \$16 \$6797 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47793 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$47794 \$153 \$6891 \$6788 \$6916 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47797 \$153 \$6827 \$6756 \$6801 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47798 \$153 \$6829 \$6789 \$6916 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47799 \$16 \$6916 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47800 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$47801 \$153 \$6872 \$6789 \$6754 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47802 \$153 \$6872 \$6756 \$6803 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47804 \$16 \$6754 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47805 \$16 \$6771 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47806 \$16 \$5932 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47807 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$47808 \$153 \$6772 \$6756 \$6805 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47809 \$153 \$6892 \$6790 \$6797 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47810 \$153 \$6671 \$5519 \$6291 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47811 \$16 \$6893 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47812 \$16 \$6797 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47813 \$16 \$6771 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47816 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$47817 \$153 \$6773 \$6756 \$6919 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47818 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$47819 \$16 \$6862 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47820 \$153 \$3199 \$5566 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$47821 \$153 \$6873 \$6906 \$6919 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47822 \$16 \$3199 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47823 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$47825 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$47827 \$153 \$6806 \$6642 \$5796 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47828 \$16 \$5796 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47829 \$16 \$5932 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47830 \$16 \$1538 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47831 \$153 \$1538 \$5702 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$47832 \$16 \$5834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47833 \$16 \$5932 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47834 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$47837 \$153 \$6874 \$5795 \$6556 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47838 \$153 \$6833 \$6698 \$5856 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47839 \$153 \$6833 \$5795 \$6616 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47841 \$16 \$5796 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47842 \$153 \$6894 \$6698 \$5796 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47845 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$47846 \$16 \$5856 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47847 \$153 \$6895 \$6585 \$5856 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47848 \$153 \$6834 \$5881 \$6617 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47849 \$153 \$6835 \$6585 \$5605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47850 \$153 \$6835 \$5625 \$6617 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47853 \$16 \$5796 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47854 \$153 \$6875 \$5625 \$6714 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47855 \$153 \$6836 \$6643 \$5796 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47856 \$153 \$6836 \$5775 \$6714 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47858 \$16 \$5605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47859 \$153 \$6837 \$6511 \$5605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47862 \$153 \$6876 \$5795 \$6558 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47863 \$153 \$6837 \$5625 \$6558 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47864 \$153 \$6838 \$6563 \$5856 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47865 \$153 \$6838 \$5795 \$6533 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47867 \$16 \$5796 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47868 \$153 \$6877 \$5795 \$6560 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47870 \$153 \$6840 \$6645 \$5796 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47872 \$153 \$6776 \$6645 \$5834 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47873 \$16 \$5834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47874 \$16 \$4837 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47875 \$16 \$5714 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47876 \$153 \$6878 \$6742 \$5714 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47880 \$16 \$5819 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47881 \$16 \$5605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47883 \$153 \$6841 \$5881 \$6715 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47884 \$16 \$5173 \$16 \$153 \$6715 VNB sky130_fd_sc_hd__inv_1
X$47885 \$153 \$6842 \$6200 \$6715 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47886 \$153 \$6843 \$6703 \$5834 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47887 \$153 \$6844 \$6200 \$6677 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47888 \$16 \$5306 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47889 \$16 \$5235 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47891 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$47892 \$16 \$1539 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47893 \$153 \$6879 \$5775 \$6677 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47894 \$153 \$1539 \$5636 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$47895 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$47896 \$16 \$5636 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47897 \$153 \$6845 \$6679 \$5636 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47899 \$153 \$6845 \$5509 \$6657 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47900 \$16 \$4834 \$16 \$153 \$6657 VNB sky130_fd_sc_hd__inv_1
X$47902 \$153 \$6896 \$6679 \$5609 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47903 \$153 \$6846 \$5635 \$6657 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47904 \$16 \$5767 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47905 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$47907 \$153 \$6880 \$5074 \$6682 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47910 \$16 \$5636 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47911 \$153 \$6848 \$6681 \$5636 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47912 \$153 \$6848 \$5509 \$6682 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47913 \$153 \$6849 \$6619 \$5786 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47915 \$153 \$6849 \$5635 \$6639 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47916 \$16 \$5786 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47918 \$153 \$6881 \$5074 \$6639 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47919 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$47920 \$16 \$5786 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47921 \$153 \$6851 \$6631 \$5786 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47922 \$153 \$6851 \$5635 \$6633 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47923 \$153 \$6852 \$6640 \$5887 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47925 \$16 \$4954 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47926 \$16 \$5609 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47927 \$153 \$6882 \$5635 \$6684 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47928 \$153 \$6897 \$6620 \$5609 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47929 \$153 \$6858 \$6620 \$5786 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47930 \$153 \$6858 \$5635 \$6565 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47933 \$16 \$5786 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47934 \$153 \$6853 \$6686 \$5786 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47935 \$153 \$6853 \$5635 \$6561 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47936 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$47937 \$16 \$5786 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47938 \$153 \$6854 \$6688 \$5786 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47939 \$16 \$5173 \$6255 \$6728 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$47940 \$16 \$5579 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47942 \$153 \$6854 \$5635 \$6601 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47943 \$16 \$5579 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47945 \$153 \$6898 \$6747 \$5718 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47946 \$16 \$5718 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47947 \$16 \$5173 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47949 \$16 \$5786 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47950 \$153 \$6899 \$6747 \$5786 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47951 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$47953 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$47954 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$47955 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$47957 \$153 \$6900 \$6859 \$7041 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47958 \$153 \$5662 \$5055 \$4579 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47960 \$153 \$5514 \$5405 \$4579 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47961 \$16 \$4579 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47962 \$16 \$4579 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47963 \$153 \$6912 \$6859 \$6979 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47964 \$16 \$6979 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47965 \$16 \$6987 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47966 \$153 \$6927 \$6781 \$6907 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47967 \$16 \$6907 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47968 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$47971 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$47972 \$153 \$6901 \$6781 \$6981 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47973 \$153 \$6901 \$6930 \$6709 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47974 \$16 \$6981 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47975 \$16 \$6988 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47977 \$153 \$6928 \$6782 \$6907 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47978 \$16 \$6907 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47979 \$16 \$7041 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47981 \$153 \$6929 \$6782 \$6979 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47982 \$153 \$6718 \$6751 \$6792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47983 \$16 \$6792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47984 \$16 \$6979 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47985 \$16 \$6989 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47987 \$153 \$6931 \$6751 \$6907 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47989 \$16 \$6907 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47990 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$47991 \$153 \$6932 \$6752 \$6907 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47992 \$153 \$6932 \$6913 \$6692 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47993 \$153 \$6900 \$6996 \$6733 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$47995 \$153 \$6933 \$6908 \$6792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$47997 \$16 \$6792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$47999 \$16 \$6909 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48000 \$153 \$6934 \$6908 \$6860 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48001 \$153 \$6884 \$6749 \$6914 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48002 \$153 \$6902 \$6785 \$6792 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48003 \$153 \$6885 \$6749 \$6795 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48006 \$16 \$6792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48007 \$16 \$6935 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48009 \$153 \$6936 \$6786 \$6907 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48010 \$16 \$6907 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48011 \$16 \$6903 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48012 \$16 \$6753 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48013 \$16 \$6910 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48014 \$153 \$6904 \$6786 \$7041 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48015 \$153 \$6904 \$6996 \$6857 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48016 \$16 \$6792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48018 \$16 \$6792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48020 \$16 \$6907 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48021 \$153 \$6937 \$6861 \$6907 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48022 \$153 \$6823 \$6794 \$6710 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48023 \$16 \$6915 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48025 \$153 \$6938 \$6796 \$6991 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48026 \$16 \$6991 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48027 \$16 \$6862 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48030 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$48032 \$153 \$6905 \$6796 \$7044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48033 \$153 \$6824 \$6906 \$6711 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48034 \$16 \$7060 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48035 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$48036 \$153 \$6650 \$6787 \$6771 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48038 \$153 \$6635 \$6787 \$6862 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48040 \$153 \$6868 \$6755 \$6771 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48041 \$153 \$6939 \$6755 \$6916 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48042 \$16 \$6771 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48043 \$16 \$6916 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48044 \$16 \$6989 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48047 \$16 \$6862 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48049 \$153 \$6917 \$6869 \$6797 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48050 \$153 \$6917 \$6906 \$6652 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48051 \$16 \$6797 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48052 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$48053 \$153 \$6940 \$6870 \$6754 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48054 \$16 \$6754 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48055 \$16 \$6771 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48058 \$153 \$6940 \$6756 \$6918 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48060 \$153 \$6941 \$6788 \$6862 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48061 \$16 \$6916 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48063 \$153 \$6828 \$6906 \$6801 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48064 \$153 \$6942 \$6789 \$6862 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48065 \$16 \$6862 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48067 \$16 \$6909 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48068 \$153 \$6802 \$6789 \$6771 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48069 \$153 \$6830 \$6906 \$6803 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48071 \$153 \$6943 \$6790 \$6916 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48072 \$153 \$6943 \$6867 \$6805 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48073 \$16 \$6916 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48077 \$16 \$6916 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48078 \$153 \$6892 \$6906 \$6805 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48079 \$153 \$6944 \$6791 \$6916 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48080 \$153 \$6944 \$6867 \$6919 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48082 \$16 \$6797 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48083 \$153 \$6873 \$6791 \$6797 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48086 \$16 \$6920 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48087 \$153 \$6832 \$6865 \$6919 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48089 \$153 \$6920 \$1538 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$48091 \$153 \$6945 \$6642 \$5605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48092 \$16 \$5605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48093 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$48095 \$153 \$6921 \$1539 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$48096 \$16 \$6921 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48097 \$153 \$6874 \$6642 \$5856 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48098 \$153 \$6946 \$6698 \$5702 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48099 \$16 \$6911 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48101 \$153 \$6911 \$1488 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$48103 \$153 \$6894 \$5775 \$6616 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48104 \$16 \$5702 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48105 \$153 \$6947 \$6585 \$5702 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48106 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$48108 \$16 \$5605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48110 \$153 \$6895 \$5795 \$6617 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48111 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$48112 \$16 \$5605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48113 \$153 \$6875 \$6643 \$5605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48115 \$16 \$5856 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48116 \$153 \$6948 \$6643 \$5856 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48117 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$48119 \$153 \$6948 \$5795 \$6714 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48120 \$16 \$5702 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48121 \$16 \$5856 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48122 \$153 \$6876 \$6511 \$5856 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48123 \$153 \$6922 \$5470 \$6558 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48124 \$16 \$5605 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48125 \$153 \$6949 \$6563 \$5605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48128 \$153 \$6949 \$5625 \$6533 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48129 \$153 \$6974 \$5470 \$6533 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48130 \$153 \$6877 \$6645 \$5856 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48131 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$48132 \$16 \$5702 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48133 \$153 \$6950 \$6645 \$5702 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48135 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$48136 \$16 \$5796 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48137 \$153 \$6951 \$6742 \$5796 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48138 \$153 \$6951 \$5775 \$6715 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48139 \$153 \$6952 \$6742 \$5605 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48140 \$16 \$5354 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48142 \$16 \$5834 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48143 \$16 \$5856 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48145 \$153 \$6953 \$6703 \$5856 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48146 \$16 \$5173 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48148 \$16 \$5796 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48149 \$153 \$6879 \$6703 \$5796 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48150 \$153 \$6954 \$6703 \$5702 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48151 \$16 \$1367 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48153 \$153 \$1367 \$5887 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$48154 \$153 \$1516 \$5609 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$48155 \$153 \$6955 \$6679 \$5963 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48157 \$153 \$6955 \$5806 \$6657 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48158 \$153 \$6956 \$6681 \$5767 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48159 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$48160 \$16 \$5963 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48161 \$153 \$6957 \$6681 \$5963 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48162 \$153 \$6957 \$5806 \$6682 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48164 \$153 \$6807 \$6619 \$5887 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48165 \$153 \$6923 \$5806 \$6639 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48167 \$16 \$5331 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48169 \$16 \$5963 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48170 \$153 \$6958 \$6631 \$5963 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48171 \$153 \$6850 \$5627 \$6633 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48173 \$153 \$6958 \$5806 \$6633 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48174 \$16 \$5963 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48176 \$16 \$6924 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48177 \$16 \$5786 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48178 \$153 \$6882 \$6640 \$5786 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48179 \$153 \$6959 \$6640 \$5609 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48180 \$16 \$5609 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48182 \$16 \$5786 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48183 \$16 \$5963 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48185 \$153 \$6960 \$6620 \$5963 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48186 \$153 \$6960 \$5806 \$6565 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48187 \$16 \$5887 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48188 \$153 \$6961 \$6686 \$5887 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48189 \$153 \$6961 \$5627 \$6561 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48190 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$48192 \$16 \$5887 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48193 \$153 \$6810 \$6688 \$5887 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48194 \$153 \$6925 \$5509 \$6601 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48195 \$153 \$6962 \$5074 \$6601 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48196 \$153 \$6926 \$5575 \$6601 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48197 \$153 \$6963 \$5806 \$6601 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48200 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$48202 \$16 \$5887 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48203 \$153 \$6964 \$6747 \$5887 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48204 \$153 \$6555 \$5509 \$6457 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48206 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$48207 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$48208 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$48209 \$153 \$2847 \$3207 \$1658 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48210 \$153 \$3091 \$3207 \$1980 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48211 \$16 \$1980 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48212 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$48213 \$153 \$3213 \$3394 \$3208 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48214 \$16 \$2024 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48217 \$153 \$3298 \$1792 \$2884 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48218 \$16 \$2180 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48220 \$16 \$1480 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48221 \$153 \$3214 \$2252 \$2884 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48222 \$16 \$1503 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48224 \$153 \$3011 \$2901 \$1687 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48225 \$16 \$1687 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48226 \$153 \$3392 \$2210 \$3056 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48227 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$48230 \$16 \$981 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48231 \$16 \$1942 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48232 \$153 \$3215 \$2252 \$3056 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48233 \$16 \$981 \$16 \$153 \$2886 VNB sky130_fd_sc_hd__inv_1
X$48235 \$153 \$3069 \$3170 \$1980 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48236 \$16 \$1980 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48238 \$16 \$1658 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48239 \$153 \$2728 \$3148 \$1980 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48241 \$16 \$1942 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48242 \$16 \$1980 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48244 \$153 \$3216 \$1943 \$3149 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48246 \$153 \$3150 \$3148 \$1658 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48247 \$16 \$1658 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48249 \$16 \$1795 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48250 \$153 \$3235 \$3093 \$1795 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48251 \$16 \$1687 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48253 \$153 \$3197 \$1815 \$3149 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48255 \$153 \$3236 \$3093 \$1658 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48256 \$16 \$3198 \$16 \$153 \$2442 VNB sky130_fd_sc_hd__clkbuf_2
X$48257 \$16 \$3198 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48259 \$153 \$3172 \$3017 \$1795 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48260 \$16 \$2006 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48261 \$16 \$1795 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48262 \$16 \$2647 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48265 \$153 \$3209 \$2064 \$3015 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48266 \$153 \$3235 \$1815 \$3015 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48267 \$16 \$1795 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48268 \$16 \$2024 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48269 \$153 \$3173 \$3071 \$1942 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48270 \$153 \$3174 \$3071 \$1687 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48271 \$16 \$1139 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48273 \$153 \$2974 \$2210 \$2889 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48274 \$153 \$3094 \$2064 \$2889 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48275 \$16 \$1815 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48276 \$153 \$153 \$2210 \$3151 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48277 \$153 \$3119 \$1943 \$2743 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48278 \$16 \$16 \$153 VNB sky130_fd_sc_hd__conb_1
X$48280 \$153 \$153 \$1815 \$3151 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48281 \$16 \$1354 \$16 \$153 \$3151 VNB sky130_fd_sc_hd__clkbuf_2
X$48284 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48285 \$153 \$3237 \$1482 \$2009 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48286 \$16 \$1496 \$2539 \$3072 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$48287 \$16 \$3096 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48288 \$153 \$3217 \$3020 \$2199 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48290 \$153 \$3217 \$2184 \$3058 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48291 \$16 \$2199 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48292 \$16 \$2539 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48296 \$153 \$3238 \$3020 \$2042 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48297 \$153 \$3238 \$1924 \$3058 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48298 \$153 \$2858 \$3005 \$1845 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48299 \$153 \$2992 \$1471 \$3058 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48300 \$16 \$1805 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48301 \$16 \$1805 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48304 \$153 \$2892 \$3144 \$1923 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48306 \$153 \$2787 \$3144 \$2199 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48307 \$16 \$2199 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48308 \$16 \$981 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48309 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$48310 \$153 \$3155 \$3006 \$1805 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48312 \$16 \$1805 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48313 \$16 \$2089 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48315 \$16 \$1965 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48317 \$153 \$3175 \$3006 \$2043 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48318 \$153 \$3175 \$1954 \$2925 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48319 \$153 \$3218 \$1924 \$2925 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48320 \$153 \$2860 \$1895 \$2327 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48321 \$16 \$1664 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48322 \$16 \$2075 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48325 \$153 \$3124 \$2026 \$2895 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48327 \$16 \$1925 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48328 \$16 \$2407 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48329 \$153 \$3157 \$2946 \$2043 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48330 \$153 \$3125 \$1806 \$2895 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48332 \$153 \$3242 \$3024 \$1923 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48334 \$16 \$1923 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48335 \$16 \$1264 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48336 \$16 \$3278 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48337 \$153 \$3176 \$3024 \$1965 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48338 \$153 \$3219 \$2026 \$3060 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48339 \$153 \$3220 \$1954 \$3060 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48340 \$153 \$3176 \$1806 \$3060 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48341 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$48343 \$16 \$2908 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48345 \$153 \$3221 \$1954 \$2908 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48347 \$153 \$3199 \$1845 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$48348 \$153 \$3200 \$2199 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$48349 \$16 \$3200 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48350 \$16 \$2199 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48351 \$16 \$3504 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48354 \$16 \$3608 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48355 \$16 \$3243 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48356 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48357 \$153 \$3178 \$1482 \$3504 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48358 \$153 \$3177 \$2184 \$2908 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48359 \$16 \$3244 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48360 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48361 \$153 \$3102 \$1482 \$3435 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48362 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48363 \$16 \$3333 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48365 \$153 \$153 \$1993 \$3061 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48366 \$153 \$153 \$1715 \$3061 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48367 \$153 \$153 \$1712 \$3061 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48369 \$16 \$3241 \$16 \$153 \$3139 VNB sky130_fd_sc_hd__clkbuf_2
X$48370 \$153 \$3127 \$3201 \$1738 \$3222 \$3103 \$1720 \$3139 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$48371 \$16 \$1578 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48374 \$153 \$3127 \$3202 \$1579 \$3223 \$3210 \$3161 \$3139 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$48375 \$16 \$1579 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48377 \$153 \$3204 \$1558 \$3203 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48378 \$153 \$3204 \$3211 \$1879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48379 \$16 \$1566 \$2935 \$3245 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$48380 \$16 \$1756 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48383 \$16 \$1585 \$16 \$153 \$3203 VNB sky130_fd_sc_hd__inv_1
X$48384 \$153 \$3275 \$3282 \$1879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48385 \$16 \$1518 \$16 \$153 \$3246 VNB sky130_fd_sc_hd__inv_1
X$48386 \$153 \$3247 \$3282 \$1969 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48388 \$153 \$3163 \$3140 \$1969 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48390 \$16 \$1647 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48391 \$16 \$3145 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48392 \$16 \$3082 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48393 \$16 \$3272 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48394 \$153 \$3224 \$1558 \$3162 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48395 \$16 \$1514 \$16 \$153 \$3162 VNB sky130_fd_sc_hd__inv_1
X$48396 \$16 \$1969 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48397 \$153 \$3179 \$3225 \$1969 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48398 \$16 \$2935 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48399 \$153 \$3225 \$1627 \$3181 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$48400 \$16 \$2105 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48402 \$153 \$3262 \$1993 \$3317 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48403 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$48404 \$153 \$3002 \$1712 \$2790 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48406 \$16 \$1969 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48407 \$153 \$3283 \$1649 \$3226 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$48408 \$153 \$3030 \$3085 \$1969 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48410 \$16 \$2098 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48411 \$153 \$3182 \$1993 \$3063 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48412 \$16 \$2935 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48413 \$16 \$1878 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48414 \$153 \$3227 \$3085 \$1878 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48415 \$153 \$3227 \$1868 \$3063 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48417 \$16 \$3248 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48418 \$16 \$1879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48419 \$16 \$1756 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48420 \$153 \$3228 \$1558 \$3296 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48422 \$153 \$3183 \$2438 \$3063 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48423 \$16 \$1228 \$16 \$153 \$3063 VNB sky130_fd_sc_hd__inv_1
X$48424 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48425 \$153 \$3161 \$1482 \$393 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48427 \$153 \$153 \$2267 \$3205 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48428 \$16 \$1378 \$16 \$153 \$3205 VNB sky130_fd_sc_hd__clkbuf_2
X$48429 \$16 \$16 \$153 VNB sky130_fd_sc_hd__conb_1
X$48430 \$153 \$153 \$2086 \$3205 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48432 \$153 \$3200 \$1973 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$48434 \$153 \$3229 \$1936 \$3186 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48435 \$153 \$3187 \$3185 \$2191 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48436 \$153 \$3187 \$2267 \$3186 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48440 \$16 \$1585 \$16 \$153 \$3167 VNB sky130_fd_sc_hd__inv_1
X$48441 \$153 \$3249 \$3212 \$2191 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48442 \$153 \$3188 \$3212 \$2031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48443 \$153 \$3250 \$1628 \$3230 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$48444 \$16 \$1566 \$2984 \$3230 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$48447 \$153 \$3189 \$2086 \$2780 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48448 \$16 \$2191 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48449 \$16 \$2984 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48451 \$16 \$1708 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48452 \$153 \$3147 \$1708 \$3190 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$48453 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$48454 \$16 \$2191 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48455 \$153 \$3191 \$3147 \$2191 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48456 \$16 \$1518 \$16 \$153 \$3192 VNB sky130_fd_sc_hd__inv_1
X$48459 \$16 \$1518 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48460 \$16 \$1647 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48461 \$153 \$3251 \$1647 \$3193 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$48463 \$16 \$2191 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48464 \$153 \$3194 \$3251 \$2191 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48465 \$16 \$1514 \$16 \$153 \$2931 VNB sky130_fd_sc_hd__inv_1
X$48466 \$153 \$3252 \$1649 \$3113 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$48469 \$153 \$3195 \$3252 \$2191 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48470 \$16 \$1121 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48471 \$153 \$3253 \$1627 \$3196 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$48472 \$153 \$3254 \$1593 \$3231 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$48474 \$153 \$3232 \$2267 \$3206 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48476 \$153 \$3233 \$2271 \$3206 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48477 \$16 \$1593 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48478 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$48480 \$153 \$3234 \$1936 \$3206 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48481 \$153 \$3115 \$2056 \$2923 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48482 \$153 \$3036 \$3090 \$2192 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48483 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$48485 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$48486 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$48487 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$48488 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$48490 \$153 \$3298 \$3207 \$1687 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48491 \$16 \$3284 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48492 \$16 \$2006 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48495 \$153 \$3285 \$1943 \$2884 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48496 \$16 \$1687 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48497 \$153 \$2937 \$3207 \$1795 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48498 \$16 \$1795 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48500 \$153 \$3286 \$3307 \$3208 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48501 \$16 \$1496 \$16 \$153 \$2884 VNB sky130_fd_sc_hd__inv_1
X$48502 \$16 \$1496 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48504 \$153 \$3268 \$3422 \$3208 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48507 \$153 \$3068 \$3170 \$1942 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48508 \$153 \$3287 \$1792 \$3056 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48509 \$16 \$1942 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48510 \$16 \$2006 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48511 \$153 \$3255 \$3170 \$2006 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48512 \$153 \$3255 \$1943 \$3056 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48515 \$153 \$3299 \$3170 \$1658 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48516 \$16 \$2006 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48517 \$153 \$3216 \$3148 \$2006 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48518 \$153 \$3301 \$3148 \$2024 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48519 \$16 \$2024 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48520 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$48522 \$153 \$3171 \$1792 \$3149 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48523 \$153 \$3209 \$3093 \$1942 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48524 \$153 \$3256 \$3093 \$2180 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48525 \$153 \$3256 \$2252 \$3015 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48526 \$16 \$2180 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48527 \$16 \$1980 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48528 \$16 \$1658 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48530 \$16 \$1264 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48531 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$48532 \$16 \$1171 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48533 \$153 \$3302 \$3017 \$1942 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48534 \$16 \$1942 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48535 \$16 \$1687 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48536 \$153 \$3303 \$3017 \$1687 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48537 \$153 \$3236 \$1547 \$3015 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48538 \$16 \$691 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48539 \$16 \$3288 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48541 \$153 \$3288 \$1795 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$48542 \$153 \$3276 \$2180 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$48543 \$16 \$3276 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48545 \$16 \$1792 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48546 \$16 \$2252 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48547 \$153 \$153 \$1792 \$3151 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48549 \$153 \$153 \$2252 \$3151 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48551 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48552 \$153 \$153 \$1943 \$3151 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48553 \$153 \$3289 \$1482 \$1815 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48554 \$16 \$1482 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48555 \$153 \$3257 \$1482 \$3540 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48558 \$153 \$3021 \$3005 \$2199 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48559 \$16 \$1496 \$16 \$153 \$3269 VNB sky130_fd_sc_hd__inv_1
X$48560 \$16 \$2199 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48561 \$16 \$1496 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48562 \$153 \$3258 \$3005 \$2089 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48563 \$153 \$3258 \$2026 \$3269 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48564 \$16 \$2089 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48565 \$16 \$2634 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48566 \$16 \$3306 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48569 \$153 \$3259 \$3005 \$1805 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48570 \$153 \$3290 \$1954 \$3269 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48572 \$153 \$3260 \$3144 \$2089 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48573 \$153 \$3259 \$1703 \$3269 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48574 \$16 \$2089 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48575 \$16 \$1923 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48578 \$153 \$3153 \$3144 \$2043 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48580 \$153 \$3154 \$3006 \$1965 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48581 \$16 \$2043 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48583 \$153 \$3218 \$3006 \$2042 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48584 \$16 \$2042 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48585 \$16 \$1751 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48587 \$153 \$3370 \$3308 \$1751 \$3305 \$3156 \$2245 \$3277 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$48588 \$16 \$2245 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48589 \$16 \$1802 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48590 \$153 \$3097 \$1895 \$2895 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48591 \$16 \$3270 \$3240 \$3309 \$162 \$16 \$153 VNB sky130_fd_sc_hd__mux2_1
X$48592 \$16 \$3310 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48593 \$16 \$3241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48594 \$153 \$3291 \$1924 \$2908 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48596 \$153 \$3370 \$3311 \$1572 \$3366 \$3278 \$2364 \$3277 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$48597 \$16 \$3366 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48598 \$16 \$2908 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48599 \$153 \$3242 \$1895 \$3060 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48600 \$153 \$3219 \$3024 \$2089 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48601 \$16 \$2089 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48602 \$16 \$1965 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48605 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$48606 \$153 \$3221 \$3077 \$2043 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48607 \$16 \$2043 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48609 \$16 \$2089 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48610 \$153 \$3158 \$3077 \$2089 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48612 \$16 \$3310 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48613 \$16 \$3241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48615 \$153 \$153 \$1895 \$3292 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48617 \$153 \$153 \$1806 \$3292 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48618 \$16 \$3199 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48619 \$16 \$2184 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48620 \$16 \$1703 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48621 \$16 \$1806 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48622 \$153 \$3243 \$2089 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$48623 \$153 \$3312 \$1482 \$1703 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48625 \$16 \$3276 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48627 \$153 \$3276 \$2098 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$48628 \$153 \$3222 \$1482 \$3079 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48629 \$153 \$153 \$1613 \$3061 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48630 \$16 \$3241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48631 \$16 \$3272 \$2820 \$3279 \$1309 \$16 \$153 VNB sky130_fd_sc_hd__mux2_1
X$48633 \$153 \$3127 \$3279 \$1578 \$3280 \$3273 \$1718 \$3139 \$16 \$16 VNB
+ sky130_fd_sc_hd__mux4_1
X$48634 \$153 \$3313 \$3281 \$1969 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48636 \$153 \$3293 \$3651 \$3160 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48637 \$153 \$3274 \$1613 \$3203 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48639 \$16 \$1543 \$2935 \$3028 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$48640 \$153 \$3274 \$3211 \$1969 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48641 \$153 \$3294 \$2092 \$3203 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48642 \$16 \$2104 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48643 \$153 \$3314 \$3282 \$2104 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48644 \$16 \$1879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48645 \$16 \$1969 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48646 \$16 \$2935 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48647 \$16 \$2098 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48649 \$153 \$3315 \$3282 \$2098 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48650 \$16 \$1969 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48651 \$16 \$2098 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48652 \$153 \$3261 \$3140 \$2098 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48653 \$153 \$3261 \$1993 \$3162 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48654 \$153 \$3486 \$1868 \$3162 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48655 \$16 \$2098 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48657 \$153 \$3262 \$3225 \$2098 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48658 \$153 \$3180 \$1613 \$2789 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48659 \$16 \$1758 \$16 \$153 \$3317 VNB sky130_fd_sc_hd__inv_1
X$48660 \$16 \$1627 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48662 \$16 \$1879 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48663 \$153 \$3318 \$3283 \$1879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48664 \$16 \$2098 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48665 \$16 \$1599 \$2935 \$3226 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$48667 \$153 \$3319 \$3283 \$2098 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48668 \$16 \$2098 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48669 \$153 \$3320 \$3322 \$2098 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48670 \$153 \$3322 \$1593 \$3321 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$48671 \$16 \$1878 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48672 \$16 \$1593 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48673 \$16 \$1475 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48676 \$153 \$3295 \$1868 \$3296 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48677 \$153 \$3297 \$1715 \$3296 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48679 \$153 \$3263 \$3085 \$1879 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48680 \$153 \$3263 \$1558 \$3063 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48681 \$16 \$1475 \$16 \$153 \$3296 VNB sky130_fd_sc_hd__inv_1
X$48682 \$153 \$153 \$1936 \$3205 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48684 \$153 \$3243 \$2191 \$16 \$16 VNB sky130_fd_sc_hd__clkbuf_16
X$48686 \$153 \$153 \$2265 \$3205 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48687 \$16 \$3243 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48688 \$16 \$1543 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48689 \$16 \$2031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48690 \$153 \$3229 \$3185 \$2031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48691 \$16 \$3200 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48692 \$16 \$1973 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48695 \$153 \$3264 \$3185 \$1973 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48696 \$153 \$3264 \$2056 \$3186 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48697 \$153 \$3166 \$3212 \$1973 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48698 \$16 \$2191 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48699 \$16 \$2031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48700 \$153 \$3249 \$2267 \$3167 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48704 \$16 \$2031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48705 \$16 \$2085 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48706 \$153 \$3323 \$3250 \$2031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48707 \$153 \$3324 \$3250 \$2085 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48708 \$153 \$3326 \$3250 \$2191 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48709 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$48712 \$16 \$2031 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48713 \$16 \$2192 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48714 \$153 \$3265 \$3147 \$2192 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48715 \$153 \$3111 \$2056 \$2920 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48716 \$153 \$3324 \$2271 \$3342 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48717 \$153 \$3191 \$2267 \$3192 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48718 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$48720 \$16 \$1973 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48722 \$153 \$2965 \$3251 \$1973 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48723 \$153 \$3168 \$2056 \$3192 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48725 \$16 \$2191 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48726 \$153 \$3266 \$3252 \$1973 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48727 \$153 \$3266 \$2056 \$3169 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48728 \$16 \$2984 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48732 \$16 \$2191 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48733 \$153 \$3232 \$3253 \$2191 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48735 \$153 \$3329 \$3254 \$2191 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48737 \$16 \$1973 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48738 \$153 \$3267 \$3253 \$1973 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48740 \$153 \$3267 \$2056 \$3206 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48741 \$16 \$2192 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48742 \$153 \$3234 \$3253 \$2031 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48743 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$48745 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$48746 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$48747 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$48748 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$48749 \$153 \$13399 \$13213 \$12294 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48750 \$16 \$12294 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48752 \$153 \$13295 \$12057 \$13336 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48753 \$16 \$12230 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48756 \$16 \$11757 \$12779 \$13367 \$16 \$153 VNB sky130_fd_sc_hd__and2_1
X$48757 \$153 \$13337 \$12134 \$13336 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48758 \$153 \$13368 \$13130 \$12236 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48759 \$153 \$13368 \$12134 \$13239 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48760 \$153 \$13338 \$11810 \$13336 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48761 \$16 \$12236 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48762 \$16 \$11898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48763 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$48766 \$153 \$13339 \$12057 \$13239 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48767 \$16 \$11898 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48768 \$153 \$13400 \$13250 \$12236 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48769 \$16 \$12294 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48770 \$153 \$13268 \$12229 \$13369 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48771 \$153 \$13296 \$12057 \$13369 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48772 \$16 \$11794 \$16 \$153 \$13369 VNB sky130_fd_sc_hd__inv_1
X$48773 \$16 \$11888 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48774 \$16 \$11794 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48776 \$16 \$11794 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48777 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$48778 \$16 \$11721 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48779 \$153 \$13370 \$13115 \$12095 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48780 \$16 \$12095 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48782 \$16 \$12230 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48783 \$153 \$13370 \$12353 \$13194 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48784 \$153 \$13340 \$12412 \$13194 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48785 \$153 \$13386 \$12412 \$13216 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48787 \$153 \$13401 \$13188 \$12294 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48788 \$16 \$12294 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48789 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$48790 \$153 \$13402 \$13272 \$12158 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48791 \$153 \$13271 \$12134 \$12926 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48792 \$16 \$12158 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48793 \$16 \$12236 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48794 \$16 \$12095 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48797 \$16 \$11485 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48798 \$153 \$13342 \$12229 \$13343 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48799 \$16 \$11485 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48800 \$153 \$13326 \$13305 \$12003 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48801 \$153 \$13158 \$12057 \$12795 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48802 \$153 \$12991 \$12134 \$12795 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48803 \$153 \$13186 \$12412 \$12795 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48805 \$16 \$11814 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48807 \$16 \$12158 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48808 \$153 \$13371 \$13298 \$12158 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48809 \$153 \$13371 \$12057 \$13345 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48810 \$153 \$13187 \$12993 \$12236 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48811 \$153 \$13387 \$12134 \$13345 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48813 \$153 \$13346 \$12229 \$13345 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48814 \$16 \$11795 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48816 \$153 \$13372 \$13347 \$12296 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48817 \$153 \$13372 \$12359 \$13373 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48818 \$16 \$11898 \$16 \$153 \$13373 VNB sky130_fd_sc_hd__inv_1
X$48819 \$153 \$13403 \$13347 \$12101 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48821 \$16 \$12101 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48822 \$16 \$12160 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48823 \$153 \$13348 \$12476 \$13105 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48824 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$48826 \$153 \$13374 \$13220 \$12296 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48827 \$16 \$12296 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48829 \$153 \$13404 \$13220 \$12044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48830 \$16 \$12044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48833 \$16 \$12101 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48834 \$16 \$11888 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48836 \$153 \$13405 \$13275 \$12296 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48837 \$16 \$11794 \$16 \$153 \$13327 VNB sky130_fd_sc_hd__inv_1
X$48839 \$153 \$13254 \$13275 \$12101 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48840 \$153 \$13388 \$12174 \$13327 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48841 \$16 \$12083 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48842 \$16 \$12101 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48843 \$16 \$12241 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48845 \$153 \$13389 \$12307 \$13240 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48846 \$16 \$12101 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48848 \$153 \$13375 \$13276 \$12044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48849 \$153 \$13375 \$12068 \$13240 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48850 \$153 \$13390 \$12363 \$13240 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48851 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$48852 \$16 \$12160 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48855 \$153 \$13328 \$13190 \$12296 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48856 \$16 \$12296 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48857 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$48858 \$153 \$13279 \$13224 \$12083 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48859 \$153 \$13349 \$12359 \$13242 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48860 \$16 \$11795 \$16 \$153 \$13242 VNB sky130_fd_sc_hd__inv_1
X$48861 \$16 \$12296 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48862 \$16 \$12083 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48863 \$16 \$11795 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48866 \$153 \$13350 \$12068 \$13242 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48867 \$16 \$12044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48869 \$16 \$11814 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48870 \$153 \$13281 \$12956 \$12160 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48871 \$153 \$13300 \$12068 \$13051 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48872 \$153 \$13377 \$13376 \$12101 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48874 \$153 \$13352 \$12476 \$13077 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48875 \$153 \$13377 \$12476 \$13243 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48876 \$16 \$12296 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48877 \$153 \$13406 \$13376 \$12296 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48878 \$153 \$13407 \$13376 \$12044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48880 \$16 \$12326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48882 \$153 \$13283 \$13330 \$12326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48883 \$153 \$13331 \$13330 \$12219 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48884 \$16 \$12219 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48885 \$16 \$11374 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48886 \$16 \$12298 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48887 \$16 \$12164 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48888 \$153 \$13391 \$13258 \$12164 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48890 \$153 \$13391 \$12217 \$13200 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48891 \$153 \$13392 \$12165 \$13244 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48892 \$16 \$12326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48893 \$153 \$13353 \$12264 \$13200 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48895 \$153 \$13408 \$13315 \$12326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48896 \$153 \$13354 \$12234 \$13245 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48899 \$16 \$12164 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48901 \$16 \$11772 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48902 \$16 \$12164 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48903 \$153 \$13393 \$12217 \$13245 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48904 \$153 \$13409 \$13316 \$12164 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48905 \$16 \$12326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48907 \$153 \$13284 \$12234 \$13302 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48908 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$48909 \$153 \$13394 \$12603 \$13302 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48912 \$16 \$12115 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48913 \$16 \$12164 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48914 \$153 \$13378 \$13285 \$12164 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48915 \$153 \$13356 \$12234 \$13203 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48916 \$153 \$13378 \$12217 \$13203 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48917 \$153 \$13357 \$12264 \$13203 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48918 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$48920 \$16 \$12326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48922 \$153 \$13038 \$13054 \$12326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48924 \$16 \$12164 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48925 \$16 \$12115 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48926 \$153 \$13286 \$13260 \$12164 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48927 \$16 \$12233 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48929 \$153 \$13359 \$12234 \$13109 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48930 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$48933 \$153 \$13287 \$12110 \$13109 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48935 \$16 \$12164 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48936 \$153 \$13410 \$13110 \$12164 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48937 \$153 \$13410 \$12217 \$13205 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48939 \$16 \$12571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48940 \$153 \$13411 \$13175 \$12571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48942 \$153 \$13261 \$13395 \$12298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48943 \$16 \$12115 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48944 \$153 \$13360 \$12217 \$13149 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48945 \$153 \$13379 \$13395 \$12115 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48946 \$153 \$13379 \$12234 \$13232 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48948 \$16 \$11983 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48951 \$16 \$11546 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48952 \$153 \$13332 \$12918 \$12010 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48953 \$16 \$12010 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48955 \$16 \$12120 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48956 \$153 \$13412 \$12918 \$12120 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48957 \$153 \$13363 \$12179 \$13362 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48958 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$48959 \$16 \$12287 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48961 \$153 \$13380 \$13094 \$12287 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48962 \$153 \$13396 \$12227 \$13056 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48963 \$153 \$13381 \$13152 \$12010 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48964 \$153 \$13380 \$12339 \$13056 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48965 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$48967 \$153 \$13397 \$12371 \$13058 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48968 \$153 \$13381 \$11942 \$13058 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48970 \$153 \$13333 \$13180 \$12384 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48972 \$16 \$12351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48973 \$16 \$12010 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48974 \$153 \$13382 \$13289 \$12010 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48977 \$153 \$13382 \$11942 \$13237 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48978 \$153 \$13263 \$13289 \$11983 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48979 \$153 \$13365 \$12182 \$13237 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48981 \$153 \$13292 \$13291 \$12010 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48982 \$16 \$12299 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48983 \$16 \$11983 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48985 \$153 \$13293 \$13291 \$11983 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48987 \$16 \$11016 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48988 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$48990 \$16 \$12299 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48991 \$153 \$13383 \$13126 \$12299 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48992 \$153 \$13383 \$12371 \$13209 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48993 \$16 \$11172 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48994 \$16 \$12299 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$48996 \$153 \$13384 \$13156 \$12299 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$48997 \$153 \$13384 \$12371 \$13248 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48998 \$153 \$13398 \$11942 \$13248 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$48999 \$16 \$11983 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49000 \$153 \$13385 \$13265 \$11983 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$49001 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$49003 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$49004 \$153 \$13366 \$11942 \$13249 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49005 \$153 \$13413 \$12119 \$13248 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49006 \$153 \$12909 \$12182 \$12980 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49007 \$153 \$13023 \$11942 \$12980 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49008 \$153 \$13021 \$12339 \$12980 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49009 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$49012 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$49013 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$49014 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$49015 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$49016 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_12
X$49019 \$153 \$13452 \$13213 \$12152 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$49020 \$16 \$12152 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49022 \$153 \$13453 \$13213 \$12095 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$49023 \$16 \$12095 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49025 \$16 \$12236 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49026 \$153 \$13414 \$13130 \$12294 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$49028 \$16 \$12294 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49030 \$153 \$13414 \$12208 \$13239 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49032 \$153 \$13415 \$13130 \$12095 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$49033 \$153 \$13415 \$12353 \$13239 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49034 \$16 \$12095 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49035 \$153 \$13456 \$13250 \$12294 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$49037 \$153 \$13434 \$12353 \$13369 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49038 \$16 \$12095 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49039 \$153 \$13416 \$13250 \$12152 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$49040 \$153 \$13416 \$12209 \$13369 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49041 \$16 \$12152 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49043 \$153 \$13417 \$13115 \$12294 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$49045 \$16 \$12294 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49046 \$153 \$13417 \$12208 \$13194 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49047 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_8
X$49048 \$153 \$13386 \$13188 \$12230 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$49049 \$153 \$13401 \$12208 \$13216 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49051 \$153 \$13435 \$12353 \$13216 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49052 \$16 \$12230 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49054 \$153 \$13458 \$13272 \$12236 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$49055 \$153 \$13341 \$12353 \$13343 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49056 \$153 \$13436 \$12209 \$13343 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49057 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$49058 \$153 \$13531 \$13305 \$12236 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$49060 \$153 \$13067 \$11810 \$12795 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49061 \$153 \$13437 \$12353 \$13215 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49062 \$153 \$13344 \$12229 \$13215 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49063 \$16 \$13215 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49064 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$49065 \$153 \$13307 \$13298 \$12003 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$49066 \$16 \$12003 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49067 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$49070 \$16 \$12095 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49071 \$153 \$13387 \$13298 \$12236 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$49072 \$16 \$12236 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49073 \$153 \$13438 \$12412 \$13345 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49074 \$16 \$11949 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49075 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$49076 \$153 \$13418 \$13347 \$12044 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$49079 \$153 \$13418 \$12068 \$13373 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49080 \$16 \$12296 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49081 \$16 \$12044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49083 \$153 \$13419 \$13347 \$12083 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$49084 \$153 \$13419 \$12174 \$13373 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49085 \$153 \$13420 \$13220 \$12241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$49088 \$153 \$13439 \$12307 \$13222 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49089 \$153 \$13420 \$12363 \$13222 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49090 \$16 \$12160 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49092 \$153 \$13404 \$12068 \$13222 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49093 \$153 \$13461 \$13275 \$12160 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$49094 \$153 \$13405 \$12359 \$13327 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49096 \$153 \$13462 \$13275 \$12241 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$49098 \$153 \$13277 \$13276 \$12101 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$49099 \$153 \$13463 \$13276 \$12295 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$49100 \$16 \$12295 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49101 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$49104 \$16 \$12044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49105 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$49107 \$153 \$13421 \$13190 \$12160 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$49108 \$153 \$13421 \$12028 \$13241 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49110 \$153 \$13165 \$12476 \$13241 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49111 \$153 \$13440 \$12307 \$13241 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49112 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$49115 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$49116 \$153 \$13441 \$12028 \$13242 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49117 \$153 \$13522 \$12155 \$13242 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49118 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$49119 \$153 \$13442 \$12363 \$13242 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49120 \$153 \$13141 \$12363 \$13049 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49121 \$16 \$12190 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49122 \$153 \$13514 \$12155 \$13051 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49124 \$153 \$13376 \$12190 \$13351 \$16 \$16 VNB sky130_fd_sc_hd__dlclkp_1
X$49125 \$153 \$13465 \$13376 \$12160 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$49126 \$153 \$13443 \$12363 \$13051 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49128 \$153 \$13329 \$13376 \$12083 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$49130 \$16 \$12083 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49131 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$49132 \$16 \$12044 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49133 \$153 \$13406 \$12359 \$13243 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49135 \$16 \$12164 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49136 \$153 \$13422 \$13330 \$12164 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$49137 \$153 \$13422 \$12217 \$13244 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49138 \$153 \$13444 \$12582 \$13244 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49141 \$153 \$13445 \$12603 \$13244 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49142 \$153 \$13423 \$13258 \$12298 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$49143 \$153 \$13423 \$12165 \$13200 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49145 \$153 \$13424 \$13258 \$12571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$49146 \$16 \$12571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49147 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$49149 \$153 \$13424 \$12309 \$13200 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49150 \$153 \$13446 \$12309 \$13245 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49151 \$153 \$13408 \$12264 \$13245 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49152 \$153 \$13393 \$13315 \$12164 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$49154 \$16 \$12571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49156 \$153 \$13515 \$12165 \$13302 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49159 \$153 \$13409 \$12217 \$13302 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49161 \$16 \$12297 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49162 \$153 \$13466 \$13316 \$12297 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$49163 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$49164 \$16 \$12571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49165 \$153 \$13468 \$13285 \$12571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$49166 \$16 \$12233 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49168 \$153 \$13469 \$13285 \$12233 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$49169 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$49170 \$16 \$12571 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49171 \$153 \$12860 \$13054 \$12571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$49172 \$153 \$13358 \$12217 \$12648 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49173 \$153 \$13447 \$12582 \$12648 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49177 \$153 \$13516 \$12165 \$13109 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49178 \$153 \$13431 \$13260 \$12233 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$49179 \$153 \$13448 \$12582 \$13109 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49181 \$16 \$12297 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49182 \$153 \$13425 \$13110 \$12297 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$49185 \$153 \$13425 \$12582 \$13205 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49186 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$49187 \$16 \$12219 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49188 \$153 \$13426 \$13395 \$12219 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$49189 \$153 \$13471 \$13395 \$12571 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$49190 \$153 \$13426 \$12110 \$13232 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49192 \$153 \$13427 \$13395 \$12326 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$49193 \$153 \$13427 \$12264 \$13232 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49194 \$16 \$12326 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49195 \$16 \$12299 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49197 \$153 \$13361 \$11881 \$13362 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49198 \$153 \$13449 \$12371 \$13362 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49200 \$16 \$11374 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49201 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$49203 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$49205 \$153 \$13412 \$12182 \$13362 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49206 \$16 \$12299 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49207 \$153 \$13474 \$13094 \$12299 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$49208 \$153 \$13432 \$13094 \$12351 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$49209 \$16 \$12351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49211 \$16 \$12299 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49213 \$153 \$13364 \$11942 \$13056 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49214 \$153 \$13397 \$13152 \$12299 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$49216 \$16 \$12299 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49217 \$153 \$13475 \$13180 \$12299 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$49218 \$153 \$13517 \$12119 \$13058 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49219 \$16 \$12384 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49221 \$153 \$13475 \$12371 \$13181 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49222 \$16 \$12198 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49223 \$16 \$12032 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49224 \$16 \$12351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49225 \$153 \$13477 \$13289 \$12351 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$49226 \$16 \$12287 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49227 \$16 \$11983 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49228 \$16 \$12120 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49229 \$153 \$13478 \$13289 \$12287 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$49230 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$49232 \$153 \$13450 \$12371 \$13237 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49233 \$16 \$12010 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49234 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
X$49235 \$153 \$13433 \$12119 \$13247 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49236 \$153 \$13428 \$13291 \$12299 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$49237 \$153 \$13428 \$12371 \$13247 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49238 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_4
X$49239 \$16 \$12303 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49240 \$16 \$12351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49242 \$153 \$13429 \$13126 \$12351 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$49243 \$153 \$13429 \$12119 \$13209 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49244 \$153 \$11868 \$10466 \$13451 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49245 \$153 \$13398 \$13156 \$12010 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$49246 \$16 \$12303 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49247 \$16 \$13451 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49248 \$16 \$12351 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49250 \$153 \$13413 \$13156 \$12351 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$49251 \$16 \$11627 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49252 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$49253 \$153 \$13385 \$11881 \$13249 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49255 \$16 \$12299 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49256 \$153 \$13430 \$13265 \$12299 \$16 \$16 VNB sky130_fd_sc_hd__dfxtp_1
X$49258 \$16 \$13451 \$16 \$153 VNB sky130_fd_sc_hd__diode_2
X$49260 \$153 \$13430 \$12371 \$13249 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49261 \$153 \$11925 \$10642 \$13451 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49262 \$153 \$11713 \$10285 \$13451 \$16 \$16 VNB sky130_fd_sc_hd__ebufn_2
X$49263 \$16 \$16 \$153 VNB sky130_fd_sc_hd__decap_6
X$49265 \$16 \$153 \$16 VNB sky130_fd_sc_hd__decap_3
.ENDS DFFRAM

.SUBCKT sky130_fd_sc_hd__mux2_1 VPB S A1 A0 X VPWR VGND VNB
M$1 \$11 S VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=76650000000P AD=158350000000P PS=785000U PD=1395000U
M$2 \$11 A0 \$8 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=76650000000P AD=193200000000P PS=785000U PD=1340000U
M$3 \$8 A1 \$12 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=193200000000P AD=44100000000P PS=1340000U PD=630000U
M$4 \$12 \$4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=44100000000P AD=69300000000P PS=630000U PD=750000U
M$5 VPWR S \$4 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=69300000000P AD=117600000000P PS=750000U PD=1400000U
M$6 X \$8 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=158350000000P PS=2520000U PD=1395000U
M$7 \$13 S VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=69300000000P
+ AD=112850000000P PS=750000U PD=1045000U
M$8 \$13 A1 \$8 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=69300000000P
+ AD=99750000000P PS=750000U PD=895000U
M$9 \$8 A0 \$14 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=99750000000P
+ AD=69300000000P PS=895000U PD=750000U
M$10 \$14 \$4 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=69300000000P AD=144900000000P PS=750000U PD=1110000U
M$11 VGND S \$4 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=144900000000P AD=109200000000P PS=1110000U PD=1360000U
M$12 X \$8 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=169000000000P AD=112850000000P PS=1820000U PD=1045000U
.ENDS sky130_fd_sc_hd__mux2_1

.SUBCKT sky130_fd_sc_hd__and2b_2 VPB A_N B VPWR VGND X VNB
M$1 \$4 A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=109200000000P AD=76650000000P PS=1360000U PD=785000U
M$2 VPWR \$4 \$7 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=76650000000P AD=60900000000P PS=785000U PD=710000U
M$3 \$7 B VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=60900000000P AD=228950000000P PS=710000U PD=1745000U
M$4 VPWR \$7 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=228950000000P AD=135000000000P PS=1745000U PD=1270000U
M$5 X \$7 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$6 VGND A_N \$4 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=109200000000P AD=109200000000P PS=1360000U PD=1360000U
M$7 \$7 \$4 \$10 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=109200000000P AD=56700000000P PS=1360000U PD=690000U
M$8 \$10 B VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=56700000000P
+ AD=101875000000P PS=690000U PD=990000U
M$9 VGND \$7 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=101875000000P
+ AD=87750000000P PS=990000U PD=920000U
M$10 X \$7 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=175500000000P PS=920000U PD=1840000U
.ENDS sky130_fd_sc_hd__and2b_2

.SUBCKT sky130_fd_sc_hd__and2_2 VPB A B VPWR X VGND VNB
M$1 VPWR A \$5 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=117600000000P AD=56700000000P PS=1400000U PD=690000U
M$2 \$5 B VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=56700000000P AD=166550000000P PS=690000U PD=1390000U
M$3 VPWR \$5 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=166550000000P AD=195000000000P PS=1390000U PD=1390000U
M$4 X \$5 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=195000000000P AD=380000000000P PS=1390000U PD=2760000U
M$5 \$5 A \$9 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=117600000000P
+ AD=56700000000P PS=1400000U PD=690000U
M$6 \$9 B VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=56700000000P
+ AD=111800000000P PS=690000U PD=1040000U
M$7 VGND \$5 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=111800000000P
+ AD=126750000000P PS=1040000U PD=1040000U
M$8 X \$5 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=126750000000P
+ AD=247000000000P PS=1040000U PD=2060000U
.ENDS sky130_fd_sc_hd__and2_2

.SUBCKT sky130_fd_sc_hd__clkbuf_4 VPB A VGND X VPWR VNB
M$1 \$3 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=265000000000P AD=165000000000P PS=2530000U PD=1330000U
M$2 VPWR \$3 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=165000000000P AD=140000000000P PS=1330000U PD=1280000U
M$3 X \$3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$4 VPWR \$3 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$5 X \$3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=300000000000P PS=1280000U PD=2600000U
M$6 \$3 A VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=111300000000P
+ AD=70350000000P PS=1370000U PD=755000U
M$7 VGND \$3 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=70350000000P
+ AD=58800000000P PS=755000U PD=700000U
M$8 X \$3 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=58800000000P PS=700000U PD=700000U
M$9 VGND \$3 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=58800000000P PS=700000U PD=700000U
M$10 X \$3 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=121800000000P PS=700000U PD=1420000U
.ENDS sky130_fd_sc_hd__clkbuf_4

.SUBCKT sky130_fd_sc_hd__and3_4 VPB A B C VGND VPWR X VNB
M$1 \$6 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=305000000000P AD=197500000000P PS=2610000U PD=1395000U
M$2 VPWR B \$6 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=197500000000P AD=140000000000P PS=1395000U PD=1280000U
M$3 \$6 C VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=177500000000P PS=1280000U PD=1355000U
M$4 VPWR \$6 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=177500000000P AD=140000000000P PS=1355000U PD=1280000U
M$5 X \$6 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$6 VPWR \$6 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$7 X \$6 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=285000000000P PS=1280000U PD=2570000U
M$8 \$6 A \$10 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=198250000000P
+ AD=128375000000P PS=1910000U PD=1045000U
M$9 \$10 B \$11 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=128375000000P AD=68250000000P PS=1045000U PD=860000U
M$10 \$11 C VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=68250000000P AD=138125000000P PS=860000U PD=1075000U
M$11 VGND \$6 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=138125000000P AD=91000000000P PS=1075000U PD=930000U
M$12 X \$6 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=91000000000P
+ AD=91000000000P PS=930000U PD=930000U
M$13 VGND \$6 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=91000000000P
+ AD=91000000000P PS=930000U PD=930000U
M$14 X \$6 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=91000000000P
+ AD=185250000000P PS=930000U PD=1870000U
.ENDS sky130_fd_sc_hd__and3_4

.SUBCKT sky130_fd_sc_hd__nor3b_4 VGND A B Y C_N VPWR VPB VNB
M$1 \$10 B \$9 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=135000000000P PS=2520000U PD=1270000U
M$2 \$9 B \$10 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$3 \$10 B \$9 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$4 \$9 B \$10 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$5 \$10 \$7 Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$6 Y \$7 \$10 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$7 \$10 \$7 Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$8 Y \$7 \$10 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$9 \$7 C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=280000000000P AD=135000000000P PS=2560000U PD=1270000U
M$10 VPWR A \$9 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$11 \$9 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$12 VPWR A \$9 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$13 \$9 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$14 \$7 C_N VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=182000000000P AD=87750000000P PS=1860000U PD=920000U
M$15 VGND A Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$16 Y A VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$17 VGND A Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$18 Y A VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=256750000000P PS=920000U PD=1440000U
M$19 VGND B Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=256750000000P
+ AD=87750000000P PS=1440000U PD=920000U
M$20 Y B VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$21 VGND B Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$22 Y B VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$23 VGND \$7 Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$24 Y \$7 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$25 VGND \$7 Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$26 Y \$7 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=169000000000P PS=920000U PD=1820000U
.ENDS sky130_fd_sc_hd__nor3b_4

.SUBCKT sky130_fd_sc_hd__and3b_4 VPB B C A_N VGND X VPWR VNB
M$1 \$10 A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=119700000000P AD=158250000000P PS=1410000U PD=1360000U
M$2 \$5 \$10 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=330000000000P AD=187500000000P PS=2660000U PD=1375000U
M$3 VPWR B \$5 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=187500000000P AD=150000000000P PS=1375000U PD=1300000U
M$4 \$5 C VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=150000000000P AD=177500000000P PS=1300000U PD=1355000U
M$5 VPWR \$5 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=177500000000P AD=145000000000P PS=1355000U PD=1290000U
M$6 X \$5 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=145000000000P AD=135000000000P PS=1290000U PD=1270000U
M$7 VPWR \$5 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=140000000000P PS=1270000U PD=1280000U
M$8 X \$5 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=158250000000P PS=1280000U PD=1360000U
M$9 \$5 \$10 \$11 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=198250000000P AD=121875000000P PS=1910000U PD=1025000U
M$10 \$11 B \$12 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=121875000000P AD=74750000000P PS=1025000U PD=880000U
M$11 \$12 C VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=74750000000P AD=138125000000P PS=880000U PD=1075000U
M$12 VGND \$5 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=138125000000P AD=91000000000P PS=1075000U PD=930000U
M$13 X \$5 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=91000000000P
+ AD=91000000000P PS=930000U PD=930000U
M$14 VGND \$5 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=91000000000P
+ AD=91000000000P PS=930000U PD=930000U
M$15 X \$5 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=91000000000P
+ AD=108375000000P PS=930000U PD=1010000U
M$16 VGND A_N \$10 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=108375000000P AD=149100000000P PS=1010000U PD=1550000U
.ENDS sky130_fd_sc_hd__and3b_4

.SUBCKT sky130_fd_sc_hd__conb_1 VPB HI|VPWR LO|VGND VNB
.ENDS sky130_fd_sc_hd__conb_1

.SUBCKT sky130_fd_sc_hd__decap_12 VPB VGND VPWR VNB
M$1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=4730000U W=870000U
+ AS=226200000000P AD=226200000000P PS=2260000U PD=2260000U
M$2 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 L=4730000U W=550000U
+ AS=143000000000P AD=143000000000P PS=1620000U PD=1620000U
.ENDS sky130_fd_sc_hd__decap_12

.SUBCKT sky130_fd_sc_hd__inv_1 VPB A VPWR VGND Y VNB
M$1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=260000000000P PS=2520000U PD=2520000U
M$2 VGND A Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=169000000000P
+ AD=169000000000P PS=1820000U PD=1820000U
.ENDS sky130_fd_sc_hd__inv_1

.SUBCKT sky130_fd_sc_hd__and4_2 VPB D C B A VPWR VGND X VNB
M$1 VPWR A \$3 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=109200000000P AD=74550000000P PS=1360000U PD=775000U
M$2 \$3 B VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=74550000000P AD=77700000000P PS=775000U PD=790000U
M$3 VPWR C \$3 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=77700000000P AD=58800000000P PS=790000U PD=700000U
M$4 \$3 D VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=58800000000P AD=279950000000P PS=700000U PD=1615000U
M$5 VPWR \$3 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=279950000000P AD=165000000000P PS=1615000U PD=1330000U
M$6 X \$3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=165000000000P AD=300000000000P PS=1330000U PD=2600000U
M$7 \$3 A \$11 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=109200000000P
+ AD=61950000000P PS=1360000U PD=715000U
M$8 \$11 B \$12 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=61950000000P
+ AD=79800000000P PS=715000U PD=800000U
M$9 \$12 C \$13 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=79800000000P
+ AD=69300000000P PS=800000U PD=750000U
M$10 \$13 D VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=69300000000P AD=175150000000P PS=750000U PD=1265000U
M$11 VGND \$3 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=175150000000P AD=107250000000P PS=1265000U PD=980000U
M$12 X \$3 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=107250000000P AD=195000000000P PS=980000U PD=1900000U
.ENDS sky130_fd_sc_hd__and4_2

.SUBCKT sky130_fd_sc_hd__mux4_1 VGND S0 X A1 A0 A3 A2 S1 VPWR VPB VNB
M$1 VPWR \$8 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=260000000000P PS=2520000U PD=2520000U
M$2 \$14 \$7 \$8 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=268800000000P AD=92087500000P PS=2120000U PD=990000U
M$3 \$13 S1 \$8 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=109200000000P AD=92087500000P PS=1360000U PD=990000U
M$4 \$21 S0 \$14 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=107900000000P AD=56700000000P PS=1360000U PD=690000U
M$5 \$14 \$12 \$24 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=56700000000P AD=90125000000P PS=690000U PD=995000U
M$6 \$24 A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=90125000000P AD=56700000000P PS=995000U PD=690000U
M$7 VPWR A2 \$21 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=56700000000P AD=109200000000P PS=690000U PD=1360000U
M$8 \$12 S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=108300000000P AD=107900000000P PS=1360000U PD=1360000U
M$9 \$19 \$12 \$13 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=109200000000P AD=56700000000P PS=1360000U PD=690000U
M$10 \$13 S0 \$20 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=56700000000P AD=107900000000P PS=690000U PD=1360000U
M$11 VPWR S1 \$7 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=109200000000P AD=109200000000P PS=1360000U PD=1360000U
M$12 \$19 A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=109200000000P AD=56700000000P PS=1360000U PD=690000U
M$13 VPWR A0 \$20 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=56700000000P AD=109200000000P PS=690000U PD=1360000U
M$14 \$14 S1 \$8 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=109200000000P AD=151025000000P PS=1360000U PD=1285000U
M$15 \$8 \$7 \$13 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=151025000000P AD=109200000000P PS=1285000U PD=1360000U
M$16 \$5 S0 \$14 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=109200000000P AD=56700000000P PS=1360000U PD=690000U
M$17 \$14 \$12 \$6 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=56700000000P AD=107950000000P PS=690000U PD=1360000U
M$18 \$5 A3 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=107900000000P AD=56700000000P PS=1360000U PD=690000U
M$19 VGND A2 \$6 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=56700000000P AD=109200000000P PS=690000U PD=1360000U
M$20 \$3 A1 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=109200000000P AD=56700000000P PS=1360000U PD=690000U
M$21 VGND A0 \$18 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=56700000000P AD=56700000000P PS=690000U PD=690000U
M$22 \$18 \$12 \$13 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=56700000000P AD=85225000000P PS=690000U PD=925000U
M$23 \$13 S0 \$3 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=85225000000P AD=109200000000P PS=925000U PD=1360000U
M$24 \$12 S0 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=109200000000P AD=109200000000P PS=1360000U PD=1360000U
M$25 VGND S1 \$7 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=109200000000P AD=109200000000P PS=1360000U PD=1360000U
M$26 VGND \$8 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=169000000000P AD=169000000000P PS=1820000U PD=1820000U
.ENDS sky130_fd_sc_hd__mux4_1

.SUBCKT sky130_fd_sc_hd__and2_1 VPB A B X VPWR VGND VNB
M$1 VPWR A \$7 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=117600000000P AD=56700000000P PS=1400000U PD=690000U
M$2 \$7 B VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=56700000000P AD=166550000000P PS=690000U PD=1390000U
M$3 VPWR \$7 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=166550000000P AD=475000000000P PS=1390000U PD=2950000U
M$4 \$7 A \$9 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=117600000000P
+ AD=56700000000P PS=1400000U PD=690000U
M$5 \$9 B VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=56700000000P
+ AD=111800000000P PS=690000U PD=1040000U
M$6 VGND \$7 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=111800000000P
+ AD=182000000000P PS=1040000U PD=1860000U
.ENDS sky130_fd_sc_hd__and2_1

.SUBCKT sky130_fd_sc_hd__dlclkp_1 VGND GCLK CLK GATE VPWR VPB VNB
M$1 \$6 \$5 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=270000000000P AD=149000000000P PS=2540000U PD=1325000U
M$2 VPWR \$6 \$7 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=640000U
+ AS=149000000000P AD=203200000000P PS=1325000U PD=1275000U
M$3 \$7 CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=640000U
+ AS=203200000000P AD=149000000000P PS=1275000U PD=1325000U
M$4 VPWR \$7 GCLK VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=149000000000P AD=260000000000P PS=1325000U PD=2520000U
M$5 \$3 CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=640000U
+ AS=166400000000P AD=86400000000P PS=1800000U PD=910000U
M$6 VPWR \$3 \$4 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=640000U
+ AS=86400000000P AD=166400000000P PS=910000U PD=1800000U
M$7 VPWR GATE \$16 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=640000U
+ AS=166400000000P AD=95750000000P PS=1800000U PD=965000U
M$8 \$16 \$4 \$5 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=95750000000P AD=98700000000P PS=965000U PD=890000U
M$9 \$5 \$3 \$17 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=98700000000P AD=44100000000P PS=890000U PD=630000U
M$10 \$17 \$6 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=44100000000P AD=109200000000P PS=630000U PD=1360000U
M$11 \$10 \$4 \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=390000U
+ AS=67125000000P AD=119200000000P PS=745000U PD=1090000U
M$12 \$10 \$6 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=67125000000P AD=118125000000P PS=745000U PD=1040000U
M$13 \$5 \$3 \$13 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=119200000000P AD=117125000000P PS=1090000U PD=1085000U
M$14 VGND \$5 \$6 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=118125000000P AD=169000000000P PS=1040000U PD=1820000U
M$15 VGND GATE \$13 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=128100000000P AD=117125000000P PS=1450000U PD=1085000U
M$16 \$7 \$6 \$9 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=109200000000P AD=44100000000P PS=1360000U PD=630000U
M$17 \$9 CLK VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=44100000000P AD=97000000000P PS=630000U PD=975000U
M$18 VGND \$7 GCLK VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=97000000000P AD=169000000000P PS=975000U PD=1820000U
M$19 \$3 CLK VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=109200000000P AD=56700000000P PS=1360000U PD=690000U
M$20 VGND \$3 \$4 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=56700000000P AD=109200000000P PS=690000U PD=1360000U
.ENDS sky130_fd_sc_hd__dlclkp_1

.SUBCKT sky130_fd_sc_hd__clkbuf_1 VPB A X VGND VPWR VNB
M$1 X \$3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=790000U
+ AS=205400000000P AD=114550000000P PS=2100000U PD=1080000U
M$2 VPWR A \$3 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=790000U
+ AS=114550000000P AD=205400000000P PS=1080000U PD=2100000U
M$3 X \$3 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=520000U AS=135200000000P
+ AD=75400000000P PS=1560000U PD=810000U
M$4 VGND A \$3 VNB sky130_fd_pr__nfet_01v8 L=150000U W=520000U AS=75400000000P
+ AD=135200000000P PS=810000U PD=1560000U
.ENDS sky130_fd_sc_hd__clkbuf_1

.SUBCKT sky130_fd_sc_hd__and4b_2 VGND B C X A_N D VPWR VPB VNB
M$1 \$3 A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=109200000000P AD=56700000000P PS=1360000U PD=690000U
M$2 VPWR \$3 \$4 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=56700000000P AD=98700000000P PS=690000U PD=890000U
M$3 \$4 B VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=98700000000P AD=128100000000P PS=890000U PD=1030000U
M$4 VPWR C \$4 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=128100000000P AD=66150000000P PS=1030000U PD=735000U
M$5 \$4 D VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=66150000000P AD=143250000000P PS=735000U PD=1330000U
M$6 VPWR \$4 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=143250000000P AD=152500000000P PS=1330000U PD=1305000U
M$7 X \$4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=152500000000P AD=260000000000P PS=1305000U PD=2520000U
M$8 \$4 \$3 \$10 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=109200000000P AD=44100000000P PS=1360000U PD=630000U
M$9 \$10 B \$9 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=44100000000P
+ AD=73500000000P PS=630000U PD=770000U
M$10 \$9 C \$8 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=73500000000P
+ AD=61950000000P PS=770000U PD=715000U
M$11 \$8 D VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=61950000000P
+ AD=103975000000P PS=715000U PD=1000000U
M$12 VGND \$4 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=103975000000P AD=99125000000P PS=1000000U PD=955000U
M$13 X \$4 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=99125000000P
+ AD=169000000000P PS=955000U PD=1820000U
M$14 VGND A_N \$3 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=109200000000P AD=109200000000P PS=1360000U PD=1360000U
.ENDS sky130_fd_sc_hd__and4b_2

.SUBCKT sky130_fd_sc_hd__and4bb_2 VGND X C D B_N A_N VPWR VPB VNB
M$1 \$3 A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=109200000000P AD=140750000000P PS=1360000U PD=1325000U
M$2 VPWR \$5 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140750000000P AD=135000000000P PS=1325000U PD=1270000U
M$3 X \$5 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=330750000000P PS=1270000U PD=1705000U
M$4 VPWR \$3 \$5 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=330750000000P AD=67200000000P PS=1705000U PD=740000U
M$5 \$5 \$13 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=67200000000P AD=58800000000P PS=740000U PD=700000U
M$6 VPWR C \$5 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=58800000000P AD=56700000000P PS=700000U PD=690000U
M$7 \$5 D VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=56700000000P AD=92400000000P PS=690000U PD=860000U
M$8 VPWR B_N \$13 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=92400000000P AD=109200000000P PS=860000U PD=1360000U
M$9 \$3 A_N VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=109200000000P AD=97000000000P PS=1360000U PD=975000U
M$10 VGND \$5 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=97000000000P
+ AD=87750000000P PS=975000U PD=920000U
M$11 X \$5 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=169000000000P PS=920000U PD=1820000U
M$12 \$5 \$3 \$11 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=109200000000P AD=44100000000P PS=1360000U PD=630000U
M$13 \$11 \$13 \$10 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=44100000000P AD=64050000000P PS=630000U PD=725000U
M$14 \$10 C \$9 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=64050000000P
+ AD=56700000000P PS=725000U PD=690000U
M$15 \$9 D VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=56700000000P
+ AD=92400000000P PS=690000U PD=860000U
M$16 VGND B_N \$13 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=92400000000P AD=109200000000P PS=860000U PD=1360000U
.ENDS sky130_fd_sc_hd__and4bb_2

.SUBCKT sky130_fd_sc_hd__nor4b_2 VGND Y A B C D_N VPWR VPB VNB
M$1 \$4 D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=109200000000P AD=109200000000P PS=1360000U PD=1360000U
M$2 \$9 C \$12 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=135000000000P PS=2520000U PD=1270000U
M$3 \$12 C \$9 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$4 \$9 \$4 Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$5 Y \$4 \$9 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$6 \$6 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=135000000000P PS=2520000U PD=1270000U
M$7 VPWR A \$6 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$8 \$6 B \$12 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$9 \$12 B \$6 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$10 \$4 D_N VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=109200000000P AD=109200000000P PS=1360000U PD=1360000U
M$11 VGND C Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=169000000000P
+ AD=87750000000P PS=1820000U PD=920000U
M$12 Y C VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$13 VGND \$4 Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$14 Y \$4 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=169000000000P PS=920000U PD=1820000U
M$15 VGND A Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=169000000000P
+ AD=87750000000P PS=1820000U PD=920000U
M$16 Y A VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$17 VGND B Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$18 Y B VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=169000000000P PS=920000U PD=1820000U
.ENDS sky130_fd_sc_hd__nor4b_2

.SUBCKT sky130_fd_sc_hd__clkbuf_2 VPB A VPWR VGND X VNB
M$1 \$6 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=265000000000P AD=162500000000P PS=2530000U PD=1325000U
M$2 VPWR \$6 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=162500000000P AD=135000000000P PS=1325000U PD=1270000U
M$3 X \$6 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$4 \$6 A VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=111300000000P
+ AD=68250000000P PS=1370000U PD=745000U
M$5 VGND \$6 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=68250000000P
+ AD=56700000000P PS=745000U PD=690000U
M$6 X \$6 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=56700000000P
+ AD=109200000000P PS=690000U PD=1360000U
.ENDS sky130_fd_sc_hd__clkbuf_2

.SUBCKT sky130_fd_sc_hd__decap_8 VPB VGND VPWR VNB
M$1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=2890000U W=870000U
+ AS=226200000000P AD=226200000000P PS=2260000U PD=2260000U
M$2 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 L=2890000U W=550000U
+ AS=143000000000P AD=143000000000P PS=1620000U PD=1620000U
.ENDS sky130_fd_sc_hd__decap_8

.SUBCKT sky130_fd_sc_hd__decap_3 VPB VGND VPWR VNB
M$1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=590000U W=870000U
+ AS=226200000000P AD=226200000000P PS=2260000U PD=2260000U
M$2 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 L=590000U W=550000U
+ AS=143000000000P AD=143000000000P PS=1620000U PD=1620000U
.ENDS sky130_fd_sc_hd__decap_3

.SUBCKT sky130_fd_sc_hd__decap_6 VPB VPWR VGND VNB
M$1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=1970000U W=870000U
+ AS=226200000000P AD=226200000000P PS=2260000U PD=2260000U
M$2 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 L=1970000U W=550000U
+ AS=143000000000P AD=143000000000P PS=1620000U PD=1620000U
.ENDS sky130_fd_sc_hd__decap_6

.SUBCKT sky130_fd_sc_hd__decap_4 VPB VGND VPWR VNB
M$1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=1050000U W=870000U
+ AS=226200000000P AD=226200000000P PS=2260000U PD=2260000U
M$2 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 L=1050000U W=550000U
+ AS=143000000000P AD=143000000000P PS=1620000U PD=1620000U
.ENDS sky130_fd_sc_hd__decap_4

.SUBCKT sky130_fd_sc_hd__diode_2 VPB DIODE VPWR VGND VNB
D$1 DIODE VNB sky130_fd_pr__diode_pw2nd_05v5 A=434700000000P P=2640000U
.ENDS sky130_fd_sc_hd__diode_2

.SUBCKT sky130_fd_sc_hd__clkbuf_16 VGND A X VPWR VPB VNB
M$1 VPWR A \$3 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=265000000000P AD=140000000000P PS=2530000U PD=1280000U
M$2 \$3 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$3 VPWR A \$3 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$4 \$3 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$5 VPWR \$3 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$6 X \$3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$7 VPWR \$3 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$8 X \$3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$9 VPWR \$3 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$10 X \$3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$11 VPWR \$3 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$12 X \$3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=137500000000P PS=1280000U PD=1275000U
M$13 VPWR \$3 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=137500000000P AD=140000000000P PS=1275000U PD=1280000U
M$14 X \$3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$15 VPWR \$3 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$16 X \$3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$17 VPWR \$3 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$18 X \$3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$19 VPWR \$3 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$20 X \$3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=265000000000P PS=1280000U PD=2530000U
M$21 VGND A \$3 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=111300000000P AD=58800000000P PS=1370000U PD=700000U
M$22 \$3 A VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=58800000000P PS=700000U PD=700000U
M$23 VGND A \$3 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=58800000000P PS=700000U PD=700000U
M$24 \$3 A VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=58800000000P PS=700000U PD=700000U
M$25 VGND \$3 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=58800000000P PS=700000U PD=700000U
M$26 X \$3 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=58800000000P PS=700000U PD=700000U
M$27 VGND \$3 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=58800000000P PS=700000U PD=700000U
M$28 X \$3 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=58800000000P PS=700000U PD=700000U
M$29 VGND \$3 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=58800000000P PS=700000U PD=700000U
M$30 X \$3 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=58800000000P PS=700000U PD=700000U
M$31 VGND \$3 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=58800000000P PS=700000U PD=700000U
M$32 X \$3 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=57750000000P PS=700000U PD=695000U
M$33 VGND \$3 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=57750000000P
+ AD=58800000000P PS=695000U PD=700000U
M$34 X \$3 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=58800000000P PS=700000U PD=700000U
M$35 VGND \$3 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=58800000000P PS=700000U PD=700000U
M$36 X \$3 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=58800000000P PS=700000U PD=700000U
M$37 VGND \$3 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=58800000000P PS=700000U PD=700000U
M$38 X \$3 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=58800000000P PS=700000U PD=700000U
M$39 VGND \$3 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=58800000000P PS=700000U PD=700000U
M$40 X \$3 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=111300000000P PS=700000U PD=1370000U
.ENDS sky130_fd_sc_hd__clkbuf_16

.SUBCKT sky130_fd_sc_hd__ebufn_2 VGND A Z TE_B VPWR VPB VNB
M$1 \$10 TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=940000U
+ AS=244400000000P AD=126900000000P PS=2400000U PD=1210000U
M$2 VPWR TE_B \$10 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=940000U
+ AS=126900000000P AD=370250000000P PS=1210000U PD=1745000U
M$3 \$10 \$3 Z VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=370250000000P AD=135000000000P PS=1745000U PD=1270000U
M$4 Z \$3 \$10 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$5 \$3 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=640000U
+ AS=166400000000P AD=120000000000P PS=1800000U PD=1015000U
M$6 VPWR TE_B \$5 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=640000U
+ AS=120000000000P AD=166400000000P PS=1015000U PD=1800000U
M$7 \$6 \$5 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=169000000000P AD=87750000000P PS=1820000U PD=920000U
M$8 VGND \$5 \$6 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=125125000000P PS=920000U PD=1035000U
M$9 \$6 \$3 Z VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=125125000000P
+ AD=87750000000P PS=1035000U PD=920000U
M$10 Z \$3 \$6 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=169000000000P PS=920000U PD=1820000U
M$11 \$3 A VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=109200000000P AD=78750000000P PS=1360000U PD=795000U
M$12 VGND TE_B \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=78750000000P AD=109200000000P PS=795000U PD=1360000U
.ENDS sky130_fd_sc_hd__ebufn_2

.SUBCKT sky130_fd_sc_hd__dfxtp_1 VGND Q CLK D VPWR VPB VNB
M$1 \$9 \$8 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=270000000000P AD=135000000000P PS=2540000U PD=1270000U
M$2 VPWR \$9 Q VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$3 VPWR D \$5 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=109200000000P AD=57750000000P PS=1360000U PD=695000U
M$4 \$5 \$4 \$6 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=57750000000P AD=68250000000P PS=695000U PD=745000U
M$5 \$6 \$3 \$17 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=68250000000P AD=76650000000P PS=745000U PD=785000U
M$6 \$17 \$7 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=76650000000P AD=178875000000P PS=785000U PD=1260000U
M$7 VPWR \$6 \$7 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=750000U
+ AS=178875000000P AD=109500000000P PS=1260000U PD=1075000U
M$8 \$7 \$3 \$8 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=109500000000P AD=56700000000P PS=1075000U PD=690000U
M$9 \$8 \$4 \$18 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=56700000000P AD=88200000000P PS=690000U PD=840000U
M$10 \$18 \$9 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=88200000000P AD=111300000000P PS=840000U PD=1370000U
M$11 \$3 CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=640000U
+ AS=166400000000P AD=86400000000P PS=1800000U PD=910000U
M$12 VPWR \$3 \$4 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=640000U
+ AS=86400000000P AD=166400000000P PS=910000U PD=1800000U
M$13 \$9 \$8 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=169000000000P AD=87750000000P PS=1820000U PD=920000U
M$14 VGND \$9 Q VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=169000000000P PS=920000U PD=1820000U
M$15 \$6 \$3 \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=360000U
+ AS=62100000000P AD=81300000000P PS=705000U PD=830000U
M$16 \$6 \$4 \$12 VNB sky130_fd_pr__nfet_01v8 L=150000U W=360000U
+ AS=62100000000P AD=69600000000P PS=705000U PD=765000U
M$17 \$8 \$4 \$7 VNB sky130_fd_pr__nfet_01v8 L=150000U W=360000U
+ AS=68400000000P AD=98900000000P PS=740000U PD=995000U
M$18 \$8 \$3 \$11 VNB sky130_fd_pr__nfet_01v8 L=150000U W=360000U
+ AS=68400000000P AD=66000000000P PS=740000U PD=745000U
M$19 VGND D \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=109200000000P AD=81300000000P PS=1360000U PD=830000U
M$20 \$12 \$7 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=69600000000P AD=120950000000P PS=765000U PD=1085000U
M$21 \$11 \$9 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=66000000000P AD=109200000000P PS=745000U PD=1360000U
M$22 VGND \$6 \$7 VNB sky130_fd_pr__nfet_01v8 L=150000U W=640000U
+ AS=120950000000P AD=98900000000P PS=1085000U PD=995000U
M$23 \$3 CLK VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=109200000000P AD=56700000000P PS=1360000U PD=690000U
M$24 VGND \$3 \$4 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=56700000000P AD=109200000000P PS=690000U PD=1360000U
.ENDS sky130_fd_sc_hd__dfxtp_1
