* Extracted by KLayout on : 15/07/2021 16:06

.SUBCKT mgmt_protect_hv
X$1 vdda1|vdda2|vssa1|vssa2|vssd mprj2_vdd_logic1 vccd
+ vdda1|vdda2|vssa1|vssa2|vssd vdda1|vdda2|vssa1|vssa2|vssd
+ vdda1|vdda2|vssa1|vssa2|vssd vdda1|vdda2|vssa1|vssa2|vssd
+ vdda1|vdda2|vssa1|vssa2|vssd vdda1|vdda2|vssa1|vssa2|vssd
+ sky130_fd_sc_hvl__lsbufhv2lv_1
X$2 vdda1|vdda2|vssa1|vssa2|vssd mprj_vdd_logic1 vccd
+ vdda1|vdda2|vssa1|vssa2|vssd vdda1|vdda2|vssa1|vssa2|vssd
+ vdda1|vdda2|vssa1|vssa2|vssd vdda1|vdda2|vssa1|vssa2|vssd
+ vdda1|vdda2|vssa1|vssa2|vssd vdda1|vdda2|vssa1|vssa2|vssd
+ sky130_fd_sc_hvl__lsbufhv2lv_1
X$3 vdda1|vdda2|vssa1|vssa2|vssd vdda1|vdda2|vssa1|vssa2|vssd
+ vdda1|vdda2|vssa1|vssa2|vssd sky130_fd_sc_hvl__conb_1
X$7 vdda1|vdda2|vssa1|vssa2|vssd vdda1|vdda2|vssa1|vssa2|vssd
+ vdda1|vdda2|vssa1|vssa2|vssd sky130_fd_sc_hvl__conb_1
.ENDS mgmt_protect_hv

.SUBCKT sky130_fd_sc_hvl__lsbufhv2lv_1 VGND X LVPWR VPWR VPB VPWR$1 A VGND$1 VNB
M$1 \$4 \$12 LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt L=150000U W=1120000U
+ AS=296800000000P AD=296800000000P PS=2770000U PD=2770000U
M$2 X \$4 LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt L=150000U W=1120000U
+ AS=296800000000P AD=156800000000P PS=2770000U PD=1400000U
M$3 LVPWR \$4 \$12 LVPWR sky130_fd_pr__pfet_01v8_hvt L=150000U W=1120000U
+ AS=156800000000P AD=296800000000P PS=1400000U PD=2770000U
M$4 VPWR$1 A \$7 VPB sky130_fd_pr__pfet_g5v0d10v5 L=500000U W=420000U
+ AS=119700000000P AD=111300000000P PS=1410000U PD=1370000U
M$5 VPWR \$7 \$3 VPB sky130_fd_pr__pfet_g5v0d10v5 L=500000U W=420000U
+ AS=119700000000P AD=111300000000P PS=1410000U PD=1370000U
M$6 X \$4 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=740000U AS=196100000000P
+ AD=196100000000P PS=2010000U PD=2010000U
M$7 \$4 \$3 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 L=500000U W=750000U
+ AS=198750000000P AD=198750000000P PS=2030000U PD=2030000U
M$8 \$12 \$7 VGND$1 VNB sky130_fd_pr__nfet_g5v0d10v5 L=500000U W=750000U
+ AS=198750000000P AD=198750000000P PS=2030000U PD=2030000U
M$9 \$4 \$3 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 L=500000U W=750000U
+ AS=198750000000P AD=198750000000P PS=2030000U PD=2030000U
M$10 \$3 \$7 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 L=500000U W=420000U
+ AS=119700000000P AD=178875000000P PS=1410000U PD=1260000U
M$11 VGND \$3 \$4 VNB sky130_fd_pr__nfet_g5v0d10v5 L=500000U W=750000U
+ AS=178875000000P AD=105000000000P PS=1260000U PD=1030000U
M$12 \$4 \$3 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 L=500000U W=750000U
+ AS=105000000000P AD=198750000000P PS=1030000U PD=2030000U
M$13 \$7 A VGND$1 VNB sky130_fd_pr__nfet_g5v0d10v5 L=500000U W=420000U
+ AS=119700000000P AD=178875000000P PS=1410000U PD=1260000U
M$14 VGND$1 \$7 \$12 VNB sky130_fd_pr__nfet_g5v0d10v5 L=500000U W=750000U
+ AS=178875000000P AD=105000000000P PS=1260000U PD=1030000U
M$15 \$12 \$7 VGND$1 VNB sky130_fd_pr__nfet_g5v0d10v5 L=500000U W=750000U
+ AS=105000000000P AD=105000000000P PS=1030000U PD=1030000U
M$16 VGND$1 \$7 \$12 VNB sky130_fd_pr__nfet_g5v0d10v5 L=500000U W=750000U
+ AS=105000000000P AD=198750000000P PS=1030000U PD=2030000U
.ENDS sky130_fd_sc_hvl__lsbufhv2lv_1

.SUBCKT sky130_fd_sc_hvl__conb_1 HI|LO|VGND|VPWR VPB VNB
R$1 HI|LO|VGND|VPWR HI|LO|VGND|VPWR 0
R$2 HI|LO|VGND|VPWR HI|LO|VGND|VPWR 0
.ENDS sky130_fd_sc_hvl__conb_1
