* Extracted by KLayout on : 15/07/2021 16:02

.SUBCKT gpio_control_block
X$1 \$2 \$1 VNB gpio_logic_high
X$2 \$3 \$57 \$2 \$55 \$4 \$4 VNB sky130_fd_sc_hd__einvp_8
X$4 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_3
X$5 \$3 \$30 \$36 \$17 \$10 \$4 \$4 VNB sky130_fd_sc_hd__dfrtp_2
X$6 \$4 \$32 \$31 \$3 \$4 VNB sky130_fd_sc_hd__buf_1
X$7 \$3 \$40 \$15 \$7 \$18 \$4 \$4 VNB sky130_fd_sc_hd__dfrtp_2
X$9 \$4 \$35 \$34 \$4 \$3 \$33 VNB sky130_fd_sc_hd__nand2b_2
X$12 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_3
X$13 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_3
X$14 \$4 \$32 \$38 \$3 \$4 VNB sky130_fd_sc_hd__buf_1
X$15 \$3 \$37 \$18 \$17 \$42 \$4 \$4 VNB sky130_fd_sc_hd__dfrtp_2
X$18 \$4 \$32 \$37 \$3 \$4 VNB sky130_fd_sc_hd__buf_1
X$20 \$3 \$41 \$35 \$7 \$21 \$4 \$4 VNB sky130_fd_sc_hd__dfstp_2
X$21 \$4 \$44 \$39 \$3 \$4 VNB sky130_fd_sc_hd__buf_1
X$23 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_3
X$24 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_4
X$25 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_3
X$27 \$3 \$11 \$8 \$7 \$10 \$4 \$4 VNB sky130_fd_sc_hd__dfrtp_2
X$29 \$3 \$12 \$13 \$7 \$24 \$4 \$4 VNB sky130_fd_sc_hd__dfrtp_2
X$30 \$4 \$4 \$3 VNB sky130_fd_sc_hd__decap_6
X$34 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_3
X$35 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_3
X$36 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_4
X$38 \$3 \$32 \$21 \$17 \$18 \$4 \$4 VNB sky130_fd_sc_hd__dfrtp_2
X$40 \$4 \$15 \$3 \$4 \$22 VNB sky130_fd_sc_hd__inv_2
X$41 \$4 \$16 \$12 \$3 \$4 VNB sky130_fd_sc_hd__buf_1
X$42 \$4 \$4 \$3 VNB sky130_fd_sc_hd__conb_1
X$43 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_8
X$45 \$4 \$14 \$4 \$3 VNB sky130_fd_sc_hd__diode_2
X$46 \$4 \$20 \$19 \$14 \$23 \$4 \$3 VNB sky130_fd_sc_hd__mux2_1
X$47 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_3
X$48 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_12
X$49 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_3
X$50 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_12
X$51 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_8
X$53 \$3 \$60 \$69 \$17 \$58 \$4 \$4 VNB sky130_fd_sc_hd__dfrtp_2
X$55 \$3 \$72 \$49 \$7 \$69 \$4 \$4 VNB sky130_fd_sc_hd__dfrtp_2
X$57 \$4 \$73 \$4 \$3 VNB sky130_fd_sc_hd__diode_2
X$58 \$4 \$70 \$23 \$73 \$71 \$4 \$3 VNB sky130_fd_sc_hd__mux2_1
X$60 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_3
X$61 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_3
X$62 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_12
X$63 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_12
X$66 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_4
X$68 \$3 \$68 \$65 \$64 \$69 \$4 \$4 VNB sky130_fd_sc_hd__dfrtp_2
X$69 \$3 \$80 \$78 \$7 \$36 \$4 \$4 VNB sky130_fd_sc_hd__dfrtp_2
X$71 \$4 \$88 \$4 \$76 \$3 VNB sky130_fd_sc_hd__dlygate4sd3_1
X$73 \$4 \$64 \$74 \$77 \$4 \$3 VNB sky130_fd_sc_hd__or2_2
X$75 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_3
X$76 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_12
X$77 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_3
X$78 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_12
X$79 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_12
X$80 \$4 \$4 \$3 VNB sky130_fd_sc_hd__decap_6
X$81 \$4 \$50 \$64 \$3 \$4 VNB sky130_fd_sc_hd__clkbuf_1
X$82 \$4 \$79 \$72 \$3 \$4 VNB sky130_fd_sc_hd__buf_1
X$83 \$4 \$79 \$80 \$3 \$4 VNB sky130_fd_sc_hd__buf_1
X$84 \$4 \$77 \$79 \$3 \$4 VNB sky130_fd_sc_hd__buf_1
X$86 \$3 \$81 \$82 \$7 \$42 \$4 \$4 VNB sky130_fd_sc_hd__dfrtp_2
X$87 \$4 \$77 \$45 \$3 \$4 VNB sky130_fd_sc_hd__buf_1
X$89 \$4 \$70 \$59 \$83 \$75 \$4 \$3 VNB sky130_fd_sc_hd__mux2_1
X$91 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_3
X$92 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_3
X$93 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_12
X$94 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_12
X$97 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_12
X$98 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_3
X$99 \$3 \$84 \$50 \$4 \$4 VNB sky130_fd_sc_hd__clkbuf_16
X$100 \$3 \$87 \$58 \$64 \$85 \$4 \$4 VNB sky130_fd_sc_hd__dfrtp_2
X$102 \$4 \$64 \$86 \$3 \$4 \$7 VNB sky130_fd_sc_hd__nor2b_2
X$103 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_3
X$104 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_12
X$105 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_3
X$106 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_12
X$109 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_12
X$110 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_12
X$111 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_4
X$113 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_8
X$115 \$4 \$62 \$3 \$4 \$57 VNB sky130_fd_sc_hd__inv_2
X$116 \$4 \$94 \$4 \$86 \$3 VNB sky130_fd_sc_hd__dlygate4sd3_1
X$117 \$4 \$76 \$4 \$94 \$3 VNB sky130_fd_sc_hd__dlygate4sd3_1
X$119 \$4 \$64 \$3 \$93 \$4 VNB sky130_fd_sc_hd__buf_2
X$121 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_3
X$122 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_12
X$123 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_3
X$124 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_8
X$125 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_3
X$126 \$4 \$50 \$17 \$3 \$4 VNB sky130_fd_sc_hd__clkbuf_1
X$129 \$4 \$45 \$54 \$3 \$4 VNB sky130_fd_sc_hd__buf_1
X$130 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_3
X$131 \$4 \$46 \$47 \$3 \$4 VNB sky130_fd_sc_hd__buf_1
X$132 \$3 \$47 \$24 \$17 \$51 \$4 \$4 VNB sky130_fd_sc_hd__dfrtp_2
X$133 \$3 \$38 \$42 \$17 \$36 \$4 \$4 VNB sky130_fd_sc_hd__dfrtp_2
X$134 \$4 \$45 \$32 \$3 \$4 VNB sky130_fd_sc_hd__buf_1
X$137 \$3 \$48 \$53 \$7 \$51 \$4 \$4 VNB sky130_fd_sc_hd__dfrtp_2
X$138 \$4 \$46 \$26 \$3 \$4 VNB sky130_fd_sc_hd__buf_1
X$139 \$4 \$44 \$40 \$3 \$4 VNB sky130_fd_sc_hd__buf_1
X$140 \$4 \$44 \$41 \$3 \$4 VNB sky130_fd_sc_hd__buf_1
X$141 \$3 \$39 \$34 \$7 \$43 \$4 \$4 VNB sky130_fd_sc_hd__dfstp_2
X$142 \$4 \$45 \$16 \$3 \$4 VNB sky130_fd_sc_hd__buf_1
X$143 \$4 \$45 \$44 \$3 \$4 VNB sky130_fd_sc_hd__buf_1
X$145 \$4 \$44 \$52 \$3 \$4 VNB sky130_fd_sc_hd__buf_1
X$147 \$4 \$44 \$48 \$3 \$4 VNB sky130_fd_sc_hd__buf_1
X$149 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_3
X$150 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_3
X$151 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_3
X$152 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_3
X$153 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_12
X$154 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_12
X$155 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_12
X$156 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_3
X$160 \$4 \$46 \$68 \$3 \$4 VNB sky130_fd_sc_hd__buf_1
X$161 \$3 \$56 \$51 \$64 \$65 \$4 \$4 VNB sky130_fd_sc_hd__dfrtp_2
X$162 \$3 \$54 \$43 \$17 \$21 \$4 \$4 VNB sky130_fd_sc_hd__dfrtp_2
X$163 \$3 \$66 \$67 \$7 \$65 \$4 \$4 VNB sky130_fd_sc_hd__dfrtp_2
X$165 \$4 \$45 \$46 \$3 \$4 VNB sky130_fd_sc_hd__buf_1
X$166 \$4 \$46 \$56 \$3 \$4 VNB sky130_fd_sc_hd__buf_1
X$167 \$4 \$46 \$60 \$3 \$4 VNB sky130_fd_sc_hd__buf_1
X$168 \$3 \$52 \$61 \$7 \$58 \$4 \$4 VNB sky130_fd_sc_hd__dfstp_2
X$169 \$3 \$62 \$5 \$63 \$4 \$4 VNB sky130_fd_sc_hd__ebufn_2
X$171 \$4 \$61 \$67 \$4 \$3 \$63 VNB sky130_fd_sc_hd__nand2b_2
X$172 \$4 \$61 \$20 \$4 \$59 \$3 VNB sky130_fd_sc_hd__and2_2
X$173 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_3
X$174 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_3
X$175 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_3
X$176 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_3
X$178 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_4
X$179 \$4 \$32 \$30 \$3 \$4 VNB sky130_fd_sc_hd__buf_1
X$180 \$3 \$26 \$28 \$17 \$24 \$4 \$4 VNB sky130_fd_sc_hd__dfrtp_2
X$181 \$3 \$31 \$10 \$17 \$28 \$4 \$4 VNB sky130_fd_sc_hd__dfrtp_2
X$182 \$3 \$27 \$25 \$7 \$28 \$4 \$4 VNB sky130_fd_sc_hd__dfrtp_2
X$184 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_12
X$185 \$4 \$4 \$3 VNB sky130_fd_sc_hd__decap_6
X$187 \$4 \$16 \$11 \$3 \$4 VNB sky130_fd_sc_hd__buf_1
X$188 \$4 \$14 \$4 \$3 VNB sky130_fd_sc_hd__diode_2
X$189 \$4 \$33 \$14 \$22 \$19 \$4 \$3 VNB sky130_fd_sc_hd__mux2_1
X$190 \$4 \$16 \$27 \$3 \$4 VNB sky130_fd_sc_hd__buf_1
X$194 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_3
X$195 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_3
X$196 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_3
X$197 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_3
X$198 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_12
X$199 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_12
X$200 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_12
X$201 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_12
X$202 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_12
X$205 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_12
X$206 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_12
X$207 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_12
X$208 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_3
X$209 \$4 \$79 \$89 \$3 \$4 VNB sky130_fd_sc_hd__buf_1
X$210 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_4
X$212 \$4 \$79 \$81 \$3 \$4 VNB sky130_fd_sc_hd__buf_1
X$214 \$4 \$16 \$87 \$3 \$4 VNB sky130_fd_sc_hd__buf_1
X$216 \$4 \$74 \$4 \$88 \$3 VNB sky130_fd_sc_hd__dlygate4sd3_1
X$217 \$4 \$91 \$4 \$3 VNB sky130_fd_sc_hd__diode_2
X$218 \$3 \$90 \$85 \$64 \$91 \$4 \$4 VNB sky130_fd_sc_hd__dfrtp_2
X$219 \$3 \$89 \$70 \$7 \$85 \$4 \$4 VNB sky130_fd_sc_hd__dfstp_2
X$221 \$4 \$74 \$3 \$92 \$4 VNB sky130_fd_sc_hd__buf_2
X$222 \$4 \$16 \$90 \$3 \$4 VNB sky130_fd_sc_hd__buf_1
X$223 \$4 \$79 \$66 \$3 \$4 VNB sky130_fd_sc_hd__buf_1
X$224 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_3
X$225 \$4 \$3 \$4 VNB sky130_fd_sc_hd__decap_3
.ENDS gpio_control_block

.SUBCKT gpio_logic_high \$1 \$2 VNB
X$1 \$1 \$2 \$1 VNB sky130_fd_sc_hd__decap_3
X$2 \$1 \$1 \$2 VNB sky130_fd_sc_hd__decap_6
X$4 \$1 \$2 \$1 VNB sky130_fd_sc_hd__decap_8
X$6 \$1 \$2 \$1 VNB sky130_fd_sc_hd__decap_3
X$7 \$1 \$2 \$1 VNB sky130_fd_sc_hd__decap_4
X$8 \$1 \$2 \$1 VNB sky130_fd_sc_hd__decap_3
X$9 \$1 \$2 \$1 VNB sky130_fd_sc_hd__decap_12
X$10 \$1 \$2 \$1 VNB sky130_fd_sc_hd__decap_3
X$11 \$1 \$1 \$2 VNB sky130_fd_sc_hd__decap_6
X$12 \$1 \$2 \$1 VNB sky130_fd_sc_hd__decap_3
X$14 \$1 \$2 \$1 VNB sky130_fd_sc_hd__decap_8
X$16 \$1 \$2 \$1 VNB sky130_fd_sc_hd__decap_3
X$17 \$1 \$2 \$1 VNB sky130_fd_sc_hd__decap_4
X$18 \$1 \$2 \$1 VNB sky130_fd_sc_hd__decap_3
X$19 \$1 \$2 \$1 VNB sky130_fd_sc_hd__decap_4
X$21 \$1 \$2 \$1 VNB sky130_fd_sc_hd__decap_3
X$22 \$1 \$2 \$1 VNB sky130_fd_sc_hd__decap_12
X$23 \$1 \$2 \$1 VNB sky130_fd_sc_hd__decap_3
X$24 \$1 \$1 \$2 VNB sky130_fd_sc_hd__decap_6
X$25 \$1 \$2 \$1 VNB sky130_fd_sc_hd__decap_3
X$27 \$1 \$2 \$1 VNB sky130_fd_sc_hd__decap_8
X$29 \$1 \$2 \$1 VNB sky130_fd_sc_hd__decap_3
X$30 \$1 \$2 \$1 VNB sky130_fd_sc_hd__decap_4
X$31 \$1 \$2 \$1 VNB sky130_fd_sc_hd__decap_3
X$33 \$1 \$1 \$2 VNB sky130_fd_sc_hd__conb_1
.ENDS gpio_logic_high

.SUBCKT sky130_fd_sc_hd__clkbuf_1 VPB A X VGND VPWR VNB
M$1 X \$3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=790000U
+ AS=205400000000P AD=114550000000P PS=2100000U PD=1080000U
M$2 VPWR A \$3 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=790000U
+ AS=114550000000P AD=205400000000P PS=1080000U PD=2100000U
M$3 X \$3 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=520000U AS=135200000000P
+ AD=75400000000P PS=1560000U PD=810000U
M$4 VGND A \$3 VNB sky130_fd_pr__nfet_01v8 L=150000U W=520000U AS=75400000000P
+ AD=135200000000P PS=810000U PD=1560000U
.ENDS sky130_fd_sc_hd__clkbuf_1

.SUBCKT sky130_fd_sc_hd__inv_2 VPB A VGND VPWR Y VNB
M$1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=135000000000P PS=2520000U PD=1270000U
M$2 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$3 VGND A Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=169000000000P
+ AD=87750000000P PS=1820000U PD=920000U
M$4 Y A VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=169000000000P PS=920000U PD=1820000U
.ENDS sky130_fd_sc_hd__inv_2

.SUBCKT sky130_fd_sc_hd__buf_2 VPB A VGND X VPWR VNB
M$1 \$3 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=640000U
+ AS=166400000000P AD=149000000000P PS=1800000U PD=1325000U
M$2 VPWR \$3 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=149000000000P AD=135000000000P PS=1325000U PD=1270000U
M$3 X \$3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=265000000000P PS=1270000U PD=2530000U
M$4 \$3 A VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=109200000000P
+ AD=97000000000P PS=1360000U PD=975000U
M$5 VGND \$3 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=97000000000P
+ AD=87750000000P PS=975000U PD=920000U
M$6 X \$3 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=172250000000P PS=920000U PD=1830000U
.ENDS sky130_fd_sc_hd__buf_2

.SUBCKT sky130_fd_sc_hd__nor2b_2 VPB B_N A VGND VPWR Y VNB
M$1 \$4 B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=109200000000P AD=109200000000P PS=1360000U PD=1360000U
M$2 \$7 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=280000000000P AD=135000000000P PS=2560000U PD=1270000U
M$3 VPWR A \$7 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$4 \$7 \$4 Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$5 Y \$4 \$7 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$6 \$4 B_N VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=109200000000P AD=109200000000P PS=1360000U PD=1360000U
M$7 VGND A Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=178750000000P
+ AD=87750000000P PS=1850000U PD=920000U
M$8 Y A VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$9 VGND \$4 Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$10 Y \$4 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=169000000000P PS=920000U PD=1820000U
.ENDS sky130_fd_sc_hd__nor2b_2

.SUBCKT sky130_fd_sc_hd__or2_2 VPB A B X VPWR VGND VNB
M$1 \$4 B \$9 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=109200000000P AD=44100000000P PS=1360000U PD=630000U
M$2 \$9 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=44100000000P AD=155750000000P PS=630000U PD=1355000U
M$3 VPWR \$4 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=155750000000P AD=135000000000P PS=1355000U PD=1270000U
M$4 X \$4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$5 VGND B \$4 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=109200000000P
+ AD=56700000000P PS=1360000U PD=690000U
M$6 \$4 A VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=56700000000P
+ AD=106750000000P PS=690000U PD=1005000U
M$7 VGND \$4 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=106750000000P
+ AD=87750000000P PS=1005000U PD=920000U
M$8 X \$4 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=169000000000P PS=920000U PD=1820000U
.ENDS sky130_fd_sc_hd__or2_2

.SUBCKT sky130_fd_sc_hd__dlygate4sd3_1 VPB A VPWR X VGND VNB
M$1 \$7 \$3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=500000U W=420000U
+ AS=109200000000P AD=140750000000P PS=1360000U PD=1325000U
M$2 VPWR \$7 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140750000000P AD=260000000000P PS=1325000U PD=2520000U
M$3 \$5 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=109200000000P AD=56700000000P PS=1360000U PD=690000U
M$4 VPWR \$5 \$3 VPB sky130_fd_pr__pfet_01v8_hvt L=500000U W=420000U
+ AS=56700000000P AD=109200000000P PS=690000U PD=1360000U
M$5 \$7 \$3 VGND VNB sky130_fd_pr__nfet_01v8 L=500000U W=420000U
+ AS=109200000000P AD=97000000000P PS=1360000U PD=975000U
M$6 VGND \$7 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=97000000000P
+ AD=169000000000P PS=975000U PD=1820000U
M$7 \$5 A VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=109200000000P
+ AD=56700000000P PS=1360000U PD=690000U
M$8 VGND \$5 \$3 VNB sky130_fd_pr__nfet_01v8 L=500000U W=420000U
+ AS=56700000000P AD=109200000000P PS=690000U PD=1360000U
.ENDS sky130_fd_sc_hd__dlygate4sd3_1

.SUBCKT sky130_fd_sc_hd__ebufn_2 VGND A Z TE_B VPWR VPB VNB
M$1 \$10 TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=940000U
+ AS=244400000000P AD=126900000000P PS=2400000U PD=1210000U
M$2 VPWR TE_B \$10 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=940000U
+ AS=126900000000P AD=370250000000P PS=1210000U PD=1745000U
M$3 \$10 \$3 Z VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=370250000000P AD=135000000000P PS=1745000U PD=1270000U
M$4 Z \$3 \$10 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$5 \$3 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=640000U
+ AS=166400000000P AD=120000000000P PS=1800000U PD=1015000U
M$6 VPWR TE_B \$5 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=640000U
+ AS=120000000000P AD=166400000000P PS=1015000U PD=1800000U
M$7 \$6 \$5 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=169000000000P AD=87750000000P PS=1820000U PD=920000U
M$8 VGND \$5 \$6 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=125125000000P PS=920000U PD=1035000U
M$9 \$6 \$3 Z VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=125125000000P
+ AD=87750000000P PS=1035000U PD=920000U
M$10 Z \$3 \$6 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=169000000000P PS=920000U PD=1820000U
M$11 \$3 A VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=109200000000P AD=78750000000P PS=1360000U PD=795000U
M$12 VGND TE_B \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=78750000000P AD=109200000000P PS=795000U PD=1360000U
.ENDS sky130_fd_sc_hd__ebufn_2

.SUBCKT sky130_fd_sc_hd__mux2_1 VPB S A1 A0 X VPWR VGND VNB
M$1 \$11 S VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=76650000000P AD=158350000000P PS=785000U PD=1395000U
M$2 \$11 A0 \$8 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=76650000000P AD=193200000000P PS=785000U PD=1340000U
M$3 \$8 A1 \$12 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=193200000000P AD=44100000000P PS=1340000U PD=630000U
M$4 \$12 \$4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=44100000000P AD=69300000000P PS=630000U PD=750000U
M$5 VPWR S \$4 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=69300000000P AD=117600000000P PS=750000U PD=1400000U
M$6 X \$8 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=158350000000P PS=2520000U PD=1395000U
M$7 \$13 S VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=69300000000P
+ AD=112850000000P PS=750000U PD=1045000U
M$8 \$13 A1 \$8 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=69300000000P
+ AD=99750000000P PS=750000U PD=895000U
M$9 \$8 A0 \$14 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=99750000000P
+ AD=69300000000P PS=895000U PD=750000U
M$10 \$14 \$4 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=69300000000P AD=144900000000P PS=750000U PD=1110000U
M$11 VGND S \$4 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=144900000000P AD=109200000000P PS=1110000U PD=1360000U
M$12 X \$8 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=169000000000P AD=112850000000P PS=1820000U PD=1045000U
.ENDS sky130_fd_sc_hd__mux2_1

.SUBCKT sky130_fd_sc_hd__diode_2 VPB DIODE VPWR VGND VNB
D$1 DIODE VNB sky130_fd_pr__diode_pw2nd_05v5 A=434700000000P P=2640000U
.ENDS sky130_fd_sc_hd__diode_2

.SUBCKT sky130_fd_sc_hd__nand2b_2 VPB B A_N VPWR VGND Y VNB
M$1 \$5 A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=109200000000P AD=146800000000P PS=1360000U PD=1340000U
M$2 VPWR \$5 Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=146800000000P AD=165000000000P PS=1340000U PD=1330000U
M$3 Y \$5 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=165000000000P AD=335000000000P PS=1330000U PD=1670000U
M$4 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=335000000000P AD=135000000000P PS=1670000U PD=1270000U
M$5 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=275000000000P PS=1270000U PD=2550000U
M$6 \$5 A_N VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=109200000000P AD=194000000000P PS=1360000U PD=1950000U
M$7 \$6 \$5 Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=169000000000P
+ AD=87750000000P PS=1820000U PD=920000U
M$8 Y \$5 \$6 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$9 \$6 B VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$10 VGND B \$6 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=169000000000P PS=920000U PD=1820000U
.ENDS sky130_fd_sc_hd__nand2b_2

.SUBCKT sky130_fd_sc_hd__clkbuf_16 VGND A X VPWR VPB VNB
M$1 VPWR A \$3 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=265000000000P AD=140000000000P PS=2530000U PD=1280000U
M$2 \$3 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$3 VPWR A \$3 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$4 \$3 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$5 VPWR \$3 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$6 X \$3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$7 VPWR \$3 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$8 X \$3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$9 VPWR \$3 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$10 X \$3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$11 VPWR \$3 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$12 X \$3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=137500000000P PS=1280000U PD=1275000U
M$13 VPWR \$3 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=137500000000P AD=140000000000P PS=1275000U PD=1280000U
M$14 X \$3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$15 VPWR \$3 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$16 X \$3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$17 VPWR \$3 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$18 X \$3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$19 VPWR \$3 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$20 X \$3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=265000000000P PS=1280000U PD=2530000U
M$21 VGND A \$3 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=111300000000P AD=58800000000P PS=1370000U PD=700000U
M$22 \$3 A VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=58800000000P PS=700000U PD=700000U
M$23 VGND A \$3 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=58800000000P PS=700000U PD=700000U
M$24 \$3 A VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=58800000000P PS=700000U PD=700000U
M$25 VGND \$3 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=58800000000P PS=700000U PD=700000U
M$26 X \$3 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=58800000000P PS=700000U PD=700000U
M$27 VGND \$3 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=58800000000P PS=700000U PD=700000U
M$28 X \$3 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=58800000000P PS=700000U PD=700000U
M$29 VGND \$3 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=58800000000P PS=700000U PD=700000U
M$30 X \$3 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=58800000000P PS=700000U PD=700000U
M$31 VGND \$3 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=58800000000P PS=700000U PD=700000U
M$32 X \$3 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=57750000000P PS=700000U PD=695000U
M$33 VGND \$3 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=57750000000P
+ AD=58800000000P PS=695000U PD=700000U
M$34 X \$3 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=58800000000P PS=700000U PD=700000U
M$35 VGND \$3 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=58800000000P PS=700000U PD=700000U
M$36 X \$3 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=58800000000P PS=700000U PD=700000U
M$37 VGND \$3 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=58800000000P PS=700000U PD=700000U
M$38 X \$3 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=58800000000P PS=700000U PD=700000U
M$39 VGND \$3 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=58800000000P PS=700000U PD=700000U
M$40 X \$3 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=111300000000P PS=700000U PD=1370000U
.ENDS sky130_fd_sc_hd__clkbuf_16

.SUBCKT sky130_fd_sc_hd__and2_2 VPB A B VPWR X VGND VNB
M$1 VPWR A \$5 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=117600000000P AD=56700000000P PS=1400000U PD=690000U
M$2 \$5 B VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=56700000000P AD=166550000000P PS=690000U PD=1390000U
M$3 VPWR \$5 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=166550000000P AD=195000000000P PS=1390000U PD=1390000U
M$4 X \$5 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=195000000000P AD=380000000000P PS=1390000U PD=2760000U
M$5 \$5 A \$9 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=117600000000P
+ AD=56700000000P PS=1400000U PD=690000U
M$6 \$9 B VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=56700000000P
+ AD=111800000000P PS=690000U PD=1040000U
M$7 VGND \$5 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=111800000000P
+ AD=126750000000P PS=1040000U PD=1040000U
M$8 X \$5 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=126750000000P
+ AD=247000000000P PS=1040000U PD=2060000U
.ENDS sky130_fd_sc_hd__and2_2

.SUBCKT sky130_fd_sc_hd__buf_1 VPB A X VGND VPWR VNB
M$1 \$3 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=790000U
+ AS=205400000000P AD=114550000000P PS=2100000U PD=1080000U
M$2 VPWR \$3 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=790000U
+ AS=114550000000P AD=205400000000P PS=1080000U PD=2100000U
M$3 \$3 A VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=520000U AS=135200000000P
+ AD=75400000000P PS=1560000U PD=810000U
M$4 VGND \$3 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=520000U AS=75400000000P
+ AD=135200000000P PS=810000U PD=1560000U
.ENDS sky130_fd_sc_hd__buf_1

.SUBCKT sky130_fd_sc_hd__dfstp_2 VGND SET_B Q CLK D VPWR VPB VNB
M$1 VPWR D \$5 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=840000U
+ AS=218400000000P AD=124950000000P PS=2200000U PD=1175000U
M$2 \$5 \$4 \$6 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=124950000000P AD=56700000000P PS=1175000U PD=690000U
M$3 \$6 \$3 \$22 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=56700000000P AD=94500000000P PS=690000U PD=870000U
M$4 \$22 \$8 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=94500000000P AD=79800000000P PS=870000U PD=800000U
M$5 VPWR SET_B \$8 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=79800000000P AD=56700000000P PS=800000U PD=690000U
M$6 \$8 \$6 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=56700000000P AD=56700000000P PS=690000U PD=690000U
M$7 VPWR \$6 \$23 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=56700000000P AD=44100000000P PS=690000U PD=630000U
M$8 \$23 \$3 \$9 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=44100000000P AD=81900000000P PS=630000U PD=810000U
M$9 \$9 \$4 \$24 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=81900000000P AD=44100000000P PS=810000U PD=630000U
M$10 \$24 \$19 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=44100000000P AD=109200000000P PS=630000U PD=1360000U
M$11 \$3 CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=640000U
+ AS=166400000000P AD=86400000000P PS=1800000U PD=910000U
M$12 VPWR \$3 \$4 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=640000U
+ AS=86400000000P AD=166400000000P PS=910000U PD=1800000U
M$13 \$10 \$9 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=135000000000P PS=2520000U PD=1270000U
M$14 VPWR \$10 Q VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$15 Q \$10 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$16 \$9 SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=109200000000P AD=120750000000P PS=1360000U PD=1165000U
M$17 VPWR \$9 \$19 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=840000U
+ AS=120750000000P AD=222600000000P PS=1165000U PD=2210000U
M$18 \$10 \$9 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=169000000000P AD=87750000000P PS=1820000U PD=920000U
M$19 VGND \$10 Q VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=87750000000P PS=920000U PD=920000U
M$20 Q \$10 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=169000000000P PS=920000U PD=1820000U
M$21 \$6 \$3 \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=360000U
+ AS=72000000000P AD=93500000000P PS=760000U PD=965000U
M$22 \$6 \$4 \$12 VNB sky130_fd_pr__nfet_01v8 L=150000U W=360000U
+ AS=72000000000P AD=67050000000P PS=760000U PD=750000U
M$23 \$12 \$8 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=67050000000P AD=88200000000P PS=750000U PD=840000U
M$24 VGND SET_B \$16 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=88200000000P AD=44100000000P PS=840000U PD=630000U
M$25 \$16 \$6 \$8 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=44100000000P AD=109200000000P PS=630000U PD=1360000U
M$26 VGND D \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=640000U
+ AS=166400000000P AD=93500000000P PS=1800000U PD=965000U
M$27 \$3 CLK VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=109200000000P AD=56700000000P PS=1360000U PD=690000U
M$28 VGND \$3 \$4 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=56700000000P AD=109200000000P PS=690000U PD=1360000U
M$29 VGND \$6 \$15 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=109200000000P AD=44100000000P PS=1360000U PD=630000U
M$30 \$15 \$4 \$9 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=44100000000P AD=73500000000P PS=630000U PD=770000U
M$31 \$9 \$3 \$13 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=73500000000P AD=44100000000P PS=770000U PD=630000U
M$32 \$13 \$19 \$14 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=44100000000P AD=44100000000P PS=630000U PD=630000U
M$33 \$14 SET_B VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=44100000000P AD=113700000000P PS=630000U PD=1010000U
M$34 VGND \$9 \$19 VNB sky130_fd_pr__nfet_01v8 L=150000U W=540000U
+ AS=113700000000P AD=140400000000P PS=1010000U PD=1600000U
.ENDS sky130_fd_sc_hd__dfstp_2

.SUBCKT sky130_fd_sc_hd__einvp_8 VGND A TE Z VPWR VPB VNB
M$1 \$8 \$5 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=940000U
+ AS=244400000000P AD=126900000000P PS=2400000U PD=1210000U
M$2 VPWR \$5 \$8 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=940000U
+ AS=126900000000P AD=126900000000P PS=1210000U PD=1210000U
M$3 \$8 \$5 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=940000U
+ AS=126900000000P AD=126900000000P PS=1210000U PD=1210000U
M$4 VPWR \$5 \$8 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=940000U
+ AS=126900000000P AD=126900000000P PS=1210000U PD=1210000U
M$5 \$8 \$5 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=940000U
+ AS=126900000000P AD=126900000000P PS=1210000U PD=1210000U
M$6 VPWR \$5 \$8 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=940000U
+ AS=126900000000P AD=126900000000P PS=1210000U PD=1210000U
M$7 \$8 \$5 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=940000U
+ AS=126900000000P AD=126900000000P PS=1210000U PD=1210000U
M$8 VPWR \$5 \$8 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=940000U
+ AS=126900000000P AD=160250000000P PS=1210000U PD=1325000U
M$9 \$8 A Z VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=160250000000P AD=135000000000P PS=1325000U PD=1270000U
M$10 Z A \$8 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$11 \$8 A Z VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$12 Z A \$8 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$13 \$8 A Z VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$14 Z A \$8 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$15 \$8 A Z VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$16 Z A \$8 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$17 \$5 TE VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=260000000000P PS=2520000U PD=2520000U
M$18 \$5 TE VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=169000000000P AD=87750000000P PS=1820000U PD=920000U
M$19 VGND TE \$6 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=94250000000P PS=920000U PD=940000U
M$20 \$6 TE VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=94250000000P AD=87750000000P PS=940000U PD=920000U
M$21 VGND TE \$6 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=87750000000P PS=920000U PD=920000U
M$22 \$6 TE VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=87750000000P PS=920000U PD=920000U
M$23 VGND TE \$6 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=87750000000P PS=920000U PD=920000U
M$24 \$6 TE VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=87750000000P PS=920000U PD=920000U
M$25 VGND TE \$6 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=87750000000P PS=920000U PD=920000U
M$26 \$6 TE VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=182000000000P PS=920000U PD=1860000U
M$27 \$6 A Z VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=169000000000P
+ AD=87750000000P PS=1820000U PD=920000U
M$28 Z A \$6 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$29 \$6 A Z VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$30 Z A \$6 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$31 \$6 A Z VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$32 Z A \$6 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$33 \$6 A Z VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$34 Z A \$6 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=182000000000P PS=920000U PD=1860000U
.ENDS sky130_fd_sc_hd__einvp_8

.SUBCKT sky130_fd_sc_hd__dfrtp_2 VGND RESET_B Q CLK D VPWR VPB VNB
M$1 VPWR D \$5 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=109200000000P AD=65100000000P PS=1360000U PD=730000U
M$2 \$5 \$4 \$6 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=65100000000P AD=72450000000P PS=730000U PD=765000U
M$3 \$6 \$3 \$19 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=72450000000P AD=115500000000P PS=765000U PD=970000U
M$4 \$19 \$17 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=115500000000P AD=70350000000P PS=970000U PD=755000U
M$5 VPWR RESET_B \$19 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=70350000000P AD=109200000000P PS=755000U PD=1360000U
M$6 VPWR \$9 Q VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=301200000000P AD=135000000000P PS=2660000U PD=1270000U
M$7 Q \$9 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$8 \$3 CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=640000U
+ AS=166400000000P AD=86400000000P PS=1800000U PD=910000U
M$9 VPWR \$3 \$4 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=640000U
+ AS=86400000000P AD=166400000000P PS=910000U PD=1800000U
M$10 VPWR \$6 \$17 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=840000U
+ AS=218400000000P AD=129150000000P PS=2200000U PD=1185000U
M$11 \$17 \$3 \$8 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=129150000000P AD=58800000000P PS=1185000U PD=700000U
M$12 \$8 \$4 \$21 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=58800000000P AD=56700000000P PS=700000U PD=690000U
M$13 \$21 \$9 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=56700000000P AD=81900000000P PS=690000U PD=810000U
M$14 VPWR RESET_B \$9 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=81900000000P AD=56700000000P PS=810000U PD=690000U
M$15 \$9 \$8 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=56700000000P AD=113400000000P PS=690000U PD=1380000U
M$16 VGND \$9 Q VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=208700000000P AD=87750000000P PS=2020000U PD=920000U
M$17 Q \$9 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=169000000000P PS=920000U PD=1820000U
M$18 \$3 CLK VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=109200000000P AD=56700000000P PS=1360000U PD=690000U
M$19 VGND \$3 \$4 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=56700000000P AD=109200000000P PS=690000U PD=1360000U
M$20 \$6 \$3 \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=360000U
+ AS=59400000000P AD=66000000000P PS=690000U PD=745000U
M$21 \$6 \$4 \$12 VNB sky130_fd_pr__nfet_01v8 L=150000U W=360000U
+ AS=59400000000P AD=140100000000P PS=690000U PD=1100000U
M$22 \$8 \$4 \$17 VNB sky130_fd_pr__nfet_01v8 L=150000U W=360000U
+ AS=71100000000P AD=99900000000P PS=755000U PD=985000U
M$23 \$8 \$3 \$13 VNB sky130_fd_pr__nfet_01v8 L=150000U W=360000U
+ AS=71100000000P AD=66900000000P PS=755000U PD=750000U
M$24 VGND D \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=220500000000P AD=66000000000P PS=1890000U PD=745000U
M$25 \$12 \$17 \$14 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=140100000000P AD=44100000000P PS=1100000U PD=630000U
M$26 \$14 RESET_B VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=44100000000P AD=134600000000P PS=630000U PD=1150000U
M$27 \$13 \$9 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=66900000000P AD=124950000000P PS=750000U PD=1015000U
M$28 VGND RESET_B \$11 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=124950000000P AD=64050000000P PS=1015000U PD=725000U
M$29 \$11 \$8 \$9 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=64050000000P AD=109200000000P PS=725000U PD=1360000U
M$30 VGND \$6 \$17 VNB sky130_fd_pr__nfet_01v8 L=150000U W=640000U
+ AS=134600000000P AD=99900000000P PS=1150000U PD=985000U
.ENDS sky130_fd_sc_hd__dfrtp_2

.SUBCKT sky130_fd_sc_hd__conb_1 VPB HI|VPWR LO|VGND VNB
R$1 LO|VGND LO|VGND 0
R$2 HI|VPWR HI|VPWR 0
.ENDS sky130_fd_sc_hd__conb_1

.SUBCKT sky130_fd_sc_hd__decap_6 VPB VPWR VGND VNB
M$1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=1970000U W=870000U
+ AS=226200000000P AD=226200000000P PS=2260000U PD=2260000U
M$2 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 L=1970000U W=550000U
+ AS=143000000000P AD=143000000000P PS=1620000U PD=1620000U
.ENDS sky130_fd_sc_hd__decap_6

.SUBCKT sky130_fd_sc_hd__decap_8 VPB VGND VPWR VNB
M$1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=2890000U W=870000U
+ AS=226200000000P AD=226200000000P PS=2260000U PD=2260000U
M$2 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 L=2890000U W=550000U
+ AS=143000000000P AD=143000000000P PS=1620000U PD=1620000U
.ENDS sky130_fd_sc_hd__decap_8

.SUBCKT sky130_fd_sc_hd__decap_4 VPB VGND VPWR VNB
M$1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=1050000U W=870000U
+ AS=226200000000P AD=226200000000P PS=2260000U PD=2260000U
M$2 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 L=1050000U W=550000U
+ AS=143000000000P AD=143000000000P PS=1620000U PD=1620000U
.ENDS sky130_fd_sc_hd__decap_4

.SUBCKT sky130_fd_sc_hd__decap_3 VPB VGND VPWR VNB
M$1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=590000U W=870000U
+ AS=226200000000P AD=226200000000P PS=2260000U PD=2260000U
M$2 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 L=590000U W=550000U
+ AS=143000000000P AD=143000000000P PS=1620000U PD=1620000U
.ENDS sky130_fd_sc_hd__decap_3

.SUBCKT sky130_fd_sc_hd__decap_12 VPB VGND VPWR VNB
M$1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=4730000U W=870000U
+ AS=226200000000P AD=226200000000P PS=2260000U PD=2260000U
M$2 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 L=4730000U W=550000U
+ AS=143000000000P AD=143000000000P PS=1620000U PD=1620000U
.ENDS sky130_fd_sc_hd__decap_12
